magic
tech sky130A
magscale 1 2
timestamp 1645353543
<< obsli1 >>
rect 552 527 224204 19601
<< obsm1 >>
rect 198 76 224204 36848
<< metal2 >>
rect 846 36688 902 37088
rect 2594 36688 2650 37088
rect 4342 36688 4398 37088
rect 6090 36688 6146 37088
rect 7838 36688 7894 37088
rect 9586 36688 9642 37088
rect 11334 36688 11390 37088
rect 13082 36688 13138 37088
rect 14830 36688 14886 37088
rect 16578 36688 16634 37088
rect 18326 36688 18382 37088
rect 20074 36688 20130 37088
rect 21914 36688 21970 37088
rect 23662 36688 23718 37088
rect 25410 36688 25466 37088
rect 27158 36688 27214 37088
rect 28906 36688 28962 37088
rect 30654 36688 30710 37088
rect 32402 36688 32458 37088
rect 34150 36688 34206 37088
rect 35898 36688 35954 37088
rect 37646 36688 37702 37088
rect 39394 36688 39450 37088
rect 41142 36688 41198 37088
rect 42982 36688 43038 37088
rect 44730 36688 44786 37088
rect 46478 36688 46534 37088
rect 48226 36688 48282 37088
rect 49974 36688 50030 37088
rect 51722 36688 51778 37088
rect 53470 36688 53526 37088
rect 55218 36688 55274 37088
rect 56966 36688 57022 37088
rect 58714 36688 58770 37088
rect 60462 36688 60518 37088
rect 62302 36688 62358 37088
rect 64050 36688 64106 37088
rect 65798 36688 65854 37088
rect 67546 36688 67602 37088
rect 69294 36688 69350 37088
rect 71042 36688 71098 37088
rect 72790 36688 72846 37088
rect 74538 36688 74594 37088
rect 76286 36688 76342 37088
rect 78034 36688 78090 37088
rect 79782 36688 79838 37088
rect 81530 36688 81586 37088
rect 83370 36688 83426 37088
rect 85118 36688 85174 37088
rect 86866 36688 86922 37088
rect 88614 36688 88670 37088
rect 90362 36688 90418 37088
rect 92110 36688 92166 37088
rect 93858 36688 93914 37088
rect 95606 36688 95662 37088
rect 97354 36688 97410 37088
rect 99102 36688 99158 37088
rect 100850 36688 100906 37088
rect 102598 36688 102654 37088
rect 104438 36688 104494 37088
rect 106186 36688 106242 37088
rect 107934 36688 107990 37088
rect 109682 36688 109738 37088
rect 111430 36688 111486 37088
rect 113178 36688 113234 37088
rect 114926 36688 114982 37088
rect 116674 36688 116730 37088
rect 118422 36688 118478 37088
rect 120170 36688 120226 37088
rect 121918 36688 121974 37088
rect 123758 36688 123814 37088
rect 125506 36688 125562 37088
rect 127254 36688 127310 37088
rect 129002 36688 129058 37088
rect 130750 36688 130806 37088
rect 132498 36688 132554 37088
rect 134246 36688 134302 37088
rect 135994 36688 136050 37088
rect 137742 36688 137798 37088
rect 139490 36688 139546 37088
rect 141238 36688 141294 37088
rect 142986 36688 143042 37088
rect 144826 36688 144882 37088
rect 146574 36688 146630 37088
rect 148322 36688 148378 37088
rect 150070 36688 150126 37088
rect 151818 36688 151874 37088
rect 153566 36688 153622 37088
rect 155314 36688 155370 37088
rect 157062 36688 157118 37088
rect 158810 36688 158866 37088
rect 160558 36688 160614 37088
rect 162306 36688 162362 37088
rect 164054 36688 164110 37088
rect 165894 36688 165950 37088
rect 167642 36688 167698 37088
rect 169390 36688 169446 37088
rect 171138 36688 171194 37088
rect 172886 36688 172942 37088
rect 174634 36688 174690 37088
rect 176382 36688 176438 37088
rect 178130 36688 178186 37088
rect 179878 36688 179934 37088
rect 181626 36688 181682 37088
rect 183374 36688 183430 37088
rect 185214 36688 185270 37088
rect 186962 36688 187018 37088
rect 188710 36688 188766 37088
rect 190458 36688 190514 37088
rect 192206 36688 192262 37088
rect 193954 36688 194010 37088
rect 195702 36688 195758 37088
rect 197450 36688 197506 37088
rect 199198 36688 199254 37088
rect 200946 36688 201002 37088
rect 202694 36688 202750 37088
rect 204442 36688 204498 37088
rect 206282 36688 206338 37088
rect 208030 36688 208086 37088
rect 209778 36688 209834 37088
rect 211526 36688 211582 37088
rect 213274 36688 213330 37088
rect 215022 36688 215078 37088
rect 216770 36688 216826 37088
rect 218518 36688 218574 37088
rect 220266 36688 220322 37088
rect 222014 36688 222070 37088
rect 223762 36688 223818 37088
rect 1766 0 1822 400
rect 5262 0 5318 400
rect 8758 0 8814 400
rect 12254 0 12310 400
rect 15750 0 15806 400
rect 19246 0 19302 400
rect 22834 0 22890 400
rect 26330 0 26386 400
rect 29826 0 29882 400
rect 33322 0 33378 400
rect 36818 0 36874 400
rect 40314 0 40370 400
rect 43902 0 43958 400
rect 47398 0 47454 400
rect 50894 0 50950 400
rect 54390 0 54446 400
rect 57886 0 57942 400
rect 61382 0 61438 400
rect 64970 0 65026 400
rect 68466 0 68522 400
rect 71962 0 72018 400
rect 75458 0 75514 400
rect 78954 0 79010 400
rect 82450 0 82506 400
rect 86038 0 86094 400
rect 89534 0 89590 400
rect 93030 0 93086 400
rect 96526 0 96582 400
rect 100022 0 100078 400
rect 103518 0 103574 400
rect 107106 0 107162 400
rect 110602 0 110658 400
rect 114098 0 114154 400
rect 117594 0 117650 400
rect 121090 0 121146 400
rect 124678 0 124734 400
rect 128174 0 128230 400
rect 131670 0 131726 400
rect 135166 0 135222 400
rect 138662 0 138718 400
rect 142158 0 142214 400
rect 145746 0 145802 400
rect 149242 0 149298 400
rect 152738 0 152794 400
rect 156234 0 156290 400
rect 159730 0 159786 400
rect 163226 0 163282 400
rect 166814 0 166870 400
rect 170310 0 170366 400
rect 173806 0 173862 400
rect 177302 0 177358 400
rect 180798 0 180854 400
rect 184294 0 184350 400
rect 187882 0 187938 400
rect 191378 0 191434 400
rect 194874 0 194930 400
rect 198370 0 198426 400
rect 201866 0 201922 400
rect 205362 0 205418 400
rect 208950 0 209006 400
rect 212446 0 212502 400
rect 215942 0 215998 400
rect 219438 0 219494 400
rect 222934 0 222990 400
<< obsm2 >>
rect 204 36632 790 36854
rect 958 36632 2538 36854
rect 2706 36632 4286 36854
rect 4454 36632 6034 36854
rect 6202 36632 7782 36854
rect 7950 36632 9530 36854
rect 9698 36632 11278 36854
rect 11446 36632 13026 36854
rect 13194 36632 14774 36854
rect 14942 36632 16522 36854
rect 16690 36632 18270 36854
rect 18438 36632 20018 36854
rect 20186 36632 21858 36854
rect 22026 36632 23606 36854
rect 23774 36632 25354 36854
rect 25522 36632 27102 36854
rect 27270 36632 28850 36854
rect 29018 36632 30598 36854
rect 30766 36632 32346 36854
rect 32514 36632 34094 36854
rect 34262 36632 35842 36854
rect 36010 36632 37590 36854
rect 37758 36632 39338 36854
rect 39506 36632 41086 36854
rect 41254 36632 42926 36854
rect 43094 36632 44674 36854
rect 44842 36632 46422 36854
rect 46590 36632 48170 36854
rect 48338 36632 49918 36854
rect 50086 36632 51666 36854
rect 51834 36632 53414 36854
rect 53582 36632 55162 36854
rect 55330 36632 56910 36854
rect 57078 36632 58658 36854
rect 58826 36632 60406 36854
rect 60574 36632 62246 36854
rect 62414 36632 63994 36854
rect 64162 36632 65742 36854
rect 65910 36632 67490 36854
rect 67658 36632 69238 36854
rect 69406 36632 70986 36854
rect 71154 36632 72734 36854
rect 72902 36632 74482 36854
rect 74650 36632 76230 36854
rect 76398 36632 77978 36854
rect 78146 36632 79726 36854
rect 79894 36632 81474 36854
rect 81642 36632 83314 36854
rect 83482 36632 85062 36854
rect 85230 36632 86810 36854
rect 86978 36632 88558 36854
rect 88726 36632 90306 36854
rect 90474 36632 92054 36854
rect 92222 36632 93802 36854
rect 93970 36632 95550 36854
rect 95718 36632 97298 36854
rect 97466 36632 99046 36854
rect 99214 36632 100794 36854
rect 100962 36632 102542 36854
rect 102710 36632 104382 36854
rect 104550 36632 106130 36854
rect 106298 36632 107878 36854
rect 108046 36632 109626 36854
rect 109794 36632 111374 36854
rect 111542 36632 113122 36854
rect 113290 36632 114870 36854
rect 115038 36632 116618 36854
rect 116786 36632 118366 36854
rect 118534 36632 120114 36854
rect 120282 36632 121862 36854
rect 122030 36632 123702 36854
rect 123870 36632 125450 36854
rect 125618 36632 127198 36854
rect 127366 36632 128946 36854
rect 129114 36632 130694 36854
rect 130862 36632 132442 36854
rect 132610 36632 134190 36854
rect 134358 36632 135938 36854
rect 136106 36632 137686 36854
rect 137854 36632 139434 36854
rect 139602 36632 141182 36854
rect 141350 36632 142930 36854
rect 143098 36632 144770 36854
rect 144938 36632 146518 36854
rect 146686 36632 148266 36854
rect 148434 36632 150014 36854
rect 150182 36632 151762 36854
rect 151930 36632 153510 36854
rect 153678 36632 155258 36854
rect 155426 36632 157006 36854
rect 157174 36632 158754 36854
rect 158922 36632 160502 36854
rect 160670 36632 162250 36854
rect 162418 36632 163998 36854
rect 164166 36632 165838 36854
rect 166006 36632 167586 36854
rect 167754 36632 169334 36854
rect 169502 36632 171082 36854
rect 171250 36632 172830 36854
rect 172998 36632 174578 36854
rect 174746 36632 176326 36854
rect 176494 36632 178074 36854
rect 178242 36632 179822 36854
rect 179990 36632 181570 36854
rect 181738 36632 183318 36854
rect 183486 36632 185158 36854
rect 185326 36632 186906 36854
rect 187074 36632 188654 36854
rect 188822 36632 190402 36854
rect 190570 36632 192150 36854
rect 192318 36632 193898 36854
rect 194066 36632 195646 36854
rect 195814 36632 197394 36854
rect 197562 36632 199142 36854
rect 199310 36632 200890 36854
rect 201058 36632 202638 36854
rect 202806 36632 204386 36854
rect 204554 36632 206226 36854
rect 206394 36632 207974 36854
rect 208142 36632 209722 36854
rect 209890 36632 211470 36854
rect 211638 36632 213218 36854
rect 213386 36632 214966 36854
rect 215134 36632 216714 36854
rect 216882 36632 218462 36854
rect 218630 36632 220210 36854
rect 220378 36632 221958 36854
rect 222126 36632 223706 36854
rect 223874 36632 224000 36854
rect 204 456 224000 36632
rect 204 31 1710 456
rect 1878 31 5206 456
rect 5374 31 8702 456
rect 8870 31 12198 456
rect 12366 31 15694 456
rect 15862 31 19190 456
rect 19358 31 22778 456
rect 22946 31 26274 456
rect 26442 31 29770 456
rect 29938 31 33266 456
rect 33434 31 36762 456
rect 36930 31 40258 456
rect 40426 31 43846 456
rect 44014 31 47342 456
rect 47510 31 50838 456
rect 51006 31 54334 456
rect 54502 31 57830 456
rect 57998 31 61326 456
rect 61494 31 64914 456
rect 65082 31 68410 456
rect 68578 31 71906 456
rect 72074 31 75402 456
rect 75570 31 78898 456
rect 79066 31 82394 456
rect 82562 31 85982 456
rect 86150 31 89478 456
rect 89646 31 92974 456
rect 93142 31 96470 456
rect 96638 31 99966 456
rect 100134 31 103462 456
rect 103630 31 107050 456
rect 107218 31 110546 456
rect 110714 31 114042 456
rect 114210 31 117538 456
rect 117706 31 121034 456
rect 121202 31 124622 456
rect 124790 31 128118 456
rect 128286 31 131614 456
rect 131782 31 135110 456
rect 135278 31 138606 456
rect 138774 31 142102 456
rect 142270 31 145690 456
rect 145858 31 149186 456
rect 149354 31 152682 456
rect 152850 31 156178 456
rect 156346 31 159674 456
rect 159842 31 163170 456
rect 163338 31 166758 456
rect 166926 31 170254 456
rect 170422 31 173750 456
rect 173918 31 177246 456
rect 177414 31 180742 456
rect 180910 31 184238 456
rect 184406 31 187826 456
rect 187994 31 191322 456
rect 191490 31 194818 456
rect 194986 31 198314 456
rect 198482 31 201810 456
rect 201978 31 205306 456
rect 205474 31 208894 456
rect 209062 31 212390 456
rect 212558 31 215886 456
rect 216054 31 219382 456
rect 219550 31 222878 456
rect 223046 31 224000 456
<< metal3 >>
rect 224356 35640 224756 35760
rect 0 34416 400 34536
rect 224356 33056 224756 33176
rect 224356 30336 224756 30456
rect 0 29112 400 29232
rect 224356 27752 224756 27872
rect 224356 25032 224756 25152
rect 0 23808 400 23928
rect 224356 22448 224756 22568
rect 224356 19728 224756 19848
rect 0 18504 400 18624
rect 224356 17144 224756 17264
rect 224356 14424 224756 14544
rect 0 13200 400 13320
rect 224356 11840 224756 11960
rect 224356 9120 224756 9240
rect 0 7896 400 8016
rect 224356 6536 224756 6656
rect 224356 3816 224756 3936
rect 0 2592 400 2712
rect 224356 1232 224756 1352
<< obsm3 >>
rect 400 35840 224356 36481
rect 400 35560 224276 35840
rect 400 34616 224356 35560
rect 480 34336 224356 34616
rect 400 33256 224356 34336
rect 400 32976 224276 33256
rect 400 30536 224356 32976
rect 400 30256 224276 30536
rect 400 29312 224356 30256
rect 480 29032 224356 29312
rect 400 27952 224356 29032
rect 400 27672 224276 27952
rect 400 25232 224356 27672
rect 400 24952 224276 25232
rect 400 24008 224356 24952
rect 480 23728 224356 24008
rect 400 22648 224356 23728
rect 400 22368 224276 22648
rect 400 19928 224356 22368
rect 400 19648 224276 19928
rect 400 18704 224356 19648
rect 480 18424 224356 18704
rect 400 17344 224356 18424
rect 400 17064 224276 17344
rect 400 14624 224356 17064
rect 400 14344 224276 14624
rect 400 13400 224356 14344
rect 480 13120 224356 13400
rect 400 12040 224356 13120
rect 400 11760 224276 12040
rect 400 9320 224356 11760
rect 400 9040 224276 9320
rect 400 8096 224356 9040
rect 480 7816 224356 8096
rect 400 6736 224356 7816
rect 400 6456 224276 6736
rect 400 4016 224356 6456
rect 400 3736 224276 4016
rect 400 2792 224356 3736
rect 480 2512 224356 2792
rect 400 1432 224356 2512
rect 400 1152 224276 1432
rect 400 35 224356 1152
<< metal4 >>
rect 1242 496 1862 36496
rect 19242 496 19862 36496
rect 37242 496 37862 36496
rect 55242 496 55862 36496
rect 73242 496 73862 36496
rect 91242 496 91862 36496
rect 109242 496 109862 36496
rect 127242 496 127862 36496
rect 145242 496 145862 36496
rect 163242 496 163862 36496
rect 181242 496 181862 36496
rect 199242 496 199862 36496
rect 217242 496 217862 36496
<< obsm4 >>
rect 3371 443 19162 35053
rect 19942 443 37162 35053
rect 37942 443 55162 35053
rect 55942 443 73162 35053
rect 73942 443 91162 35053
rect 91942 443 109162 35053
rect 109942 443 127162 35053
rect 127942 443 145162 35053
rect 145942 443 163162 35053
rect 163942 443 181162 35053
rect 181942 443 199162 35053
rect 199942 443 215405 35053
<< labels >>
rlabel metal3 s 224356 25032 224756 25152 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 224356 27752 224756 27872 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 224356 30336 224756 30456 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 224356 33056 224756 33176 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 224356 35640 224756 35760 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 0 7896 400 8016 6 A1[0]
port 6 nsew signal input
rlabel metal3 s 0 13200 400 13320 6 A1[1]
port 7 nsew signal input
rlabel metal3 s 0 18504 400 18624 6 A1[2]
port 8 nsew signal input
rlabel metal3 s 0 23808 400 23928 6 A1[3]
port 9 nsew signal input
rlabel metal3 s 0 29112 400 29232 6 A1[4]
port 10 nsew signal input
rlabel metal3 s 0 2592 400 2712 6 CLK
port 11 nsew signal input
rlabel metal2 s 1766 0 1822 400 6 Di0[0]
port 12 nsew signal input
rlabel metal2 s 36818 0 36874 400 6 Di0[10]
port 13 nsew signal input
rlabel metal2 s 40314 0 40370 400 6 Di0[11]
port 14 nsew signal input
rlabel metal2 s 43902 0 43958 400 6 Di0[12]
port 15 nsew signal input
rlabel metal2 s 47398 0 47454 400 6 Di0[13]
port 16 nsew signal input
rlabel metal2 s 50894 0 50950 400 6 Di0[14]
port 17 nsew signal input
rlabel metal2 s 54390 0 54446 400 6 Di0[15]
port 18 nsew signal input
rlabel metal2 s 57886 0 57942 400 6 Di0[16]
port 19 nsew signal input
rlabel metal2 s 61382 0 61438 400 6 Di0[17]
port 20 nsew signal input
rlabel metal2 s 64970 0 65026 400 6 Di0[18]
port 21 nsew signal input
rlabel metal2 s 68466 0 68522 400 6 Di0[19]
port 22 nsew signal input
rlabel metal2 s 5262 0 5318 400 6 Di0[1]
port 23 nsew signal input
rlabel metal2 s 71962 0 72018 400 6 Di0[20]
port 24 nsew signal input
rlabel metal2 s 75458 0 75514 400 6 Di0[21]
port 25 nsew signal input
rlabel metal2 s 78954 0 79010 400 6 Di0[22]
port 26 nsew signal input
rlabel metal2 s 82450 0 82506 400 6 Di0[23]
port 27 nsew signal input
rlabel metal2 s 86038 0 86094 400 6 Di0[24]
port 28 nsew signal input
rlabel metal2 s 89534 0 89590 400 6 Di0[25]
port 29 nsew signal input
rlabel metal2 s 93030 0 93086 400 6 Di0[26]
port 30 nsew signal input
rlabel metal2 s 96526 0 96582 400 6 Di0[27]
port 31 nsew signal input
rlabel metal2 s 100022 0 100078 400 6 Di0[28]
port 32 nsew signal input
rlabel metal2 s 103518 0 103574 400 6 Di0[29]
port 33 nsew signal input
rlabel metal2 s 8758 0 8814 400 6 Di0[2]
port 34 nsew signal input
rlabel metal2 s 107106 0 107162 400 6 Di0[30]
port 35 nsew signal input
rlabel metal2 s 110602 0 110658 400 6 Di0[31]
port 36 nsew signal input
rlabel metal2 s 114098 0 114154 400 6 Di0[32]
port 37 nsew signal input
rlabel metal2 s 117594 0 117650 400 6 Di0[33]
port 38 nsew signal input
rlabel metal2 s 121090 0 121146 400 6 Di0[34]
port 39 nsew signal input
rlabel metal2 s 124678 0 124734 400 6 Di0[35]
port 40 nsew signal input
rlabel metal2 s 128174 0 128230 400 6 Di0[36]
port 41 nsew signal input
rlabel metal2 s 131670 0 131726 400 6 Di0[37]
port 42 nsew signal input
rlabel metal2 s 135166 0 135222 400 6 Di0[38]
port 43 nsew signal input
rlabel metal2 s 138662 0 138718 400 6 Di0[39]
port 44 nsew signal input
rlabel metal2 s 12254 0 12310 400 6 Di0[3]
port 45 nsew signal input
rlabel metal2 s 142158 0 142214 400 6 Di0[40]
port 46 nsew signal input
rlabel metal2 s 145746 0 145802 400 6 Di0[41]
port 47 nsew signal input
rlabel metal2 s 149242 0 149298 400 6 Di0[42]
port 48 nsew signal input
rlabel metal2 s 152738 0 152794 400 6 Di0[43]
port 49 nsew signal input
rlabel metal2 s 156234 0 156290 400 6 Di0[44]
port 50 nsew signal input
rlabel metal2 s 159730 0 159786 400 6 Di0[45]
port 51 nsew signal input
rlabel metal2 s 163226 0 163282 400 6 Di0[46]
port 52 nsew signal input
rlabel metal2 s 166814 0 166870 400 6 Di0[47]
port 53 nsew signal input
rlabel metal2 s 170310 0 170366 400 6 Di0[48]
port 54 nsew signal input
rlabel metal2 s 173806 0 173862 400 6 Di0[49]
port 55 nsew signal input
rlabel metal2 s 15750 0 15806 400 6 Di0[4]
port 56 nsew signal input
rlabel metal2 s 177302 0 177358 400 6 Di0[50]
port 57 nsew signal input
rlabel metal2 s 180798 0 180854 400 6 Di0[51]
port 58 nsew signal input
rlabel metal2 s 184294 0 184350 400 6 Di0[52]
port 59 nsew signal input
rlabel metal2 s 187882 0 187938 400 6 Di0[53]
port 60 nsew signal input
rlabel metal2 s 191378 0 191434 400 6 Di0[54]
port 61 nsew signal input
rlabel metal2 s 194874 0 194930 400 6 Di0[55]
port 62 nsew signal input
rlabel metal2 s 198370 0 198426 400 6 Di0[56]
port 63 nsew signal input
rlabel metal2 s 201866 0 201922 400 6 Di0[57]
port 64 nsew signal input
rlabel metal2 s 205362 0 205418 400 6 Di0[58]
port 65 nsew signal input
rlabel metal2 s 208950 0 209006 400 6 Di0[59]
port 66 nsew signal input
rlabel metal2 s 19246 0 19302 400 6 Di0[5]
port 67 nsew signal input
rlabel metal2 s 212446 0 212502 400 6 Di0[60]
port 68 nsew signal input
rlabel metal2 s 215942 0 215998 400 6 Di0[61]
port 69 nsew signal input
rlabel metal2 s 219438 0 219494 400 6 Di0[62]
port 70 nsew signal input
rlabel metal2 s 222934 0 222990 400 6 Di0[63]
port 71 nsew signal input
rlabel metal2 s 22834 0 22890 400 6 Di0[6]
port 72 nsew signal input
rlabel metal2 s 26330 0 26386 400 6 Di0[7]
port 73 nsew signal input
rlabel metal2 s 29826 0 29882 400 6 Di0[8]
port 74 nsew signal input
rlabel metal2 s 33322 0 33378 400 6 Di0[9]
port 75 nsew signal input
rlabel metal2 s 846 36688 902 37088 6 Do0[0]
port 76 nsew signal output
rlabel metal2 s 18326 36688 18382 37088 6 Do0[10]
port 77 nsew signal output
rlabel metal2 s 21914 36688 21970 37088 6 Do0[11]
port 78 nsew signal output
rlabel metal2 s 25410 36688 25466 37088 6 Do0[12]
port 79 nsew signal output
rlabel metal2 s 28906 36688 28962 37088 6 Do0[13]
port 80 nsew signal output
rlabel metal2 s 32402 36688 32458 37088 6 Do0[14]
port 81 nsew signal output
rlabel metal2 s 35898 36688 35954 37088 6 Do0[15]
port 82 nsew signal output
rlabel metal2 s 39394 36688 39450 37088 6 Do0[16]
port 83 nsew signal output
rlabel metal2 s 42982 36688 43038 37088 6 Do0[17]
port 84 nsew signal output
rlabel metal2 s 46478 36688 46534 37088 6 Do0[18]
port 85 nsew signal output
rlabel metal2 s 49974 36688 50030 37088 6 Do0[19]
port 86 nsew signal output
rlabel metal2 s 2594 36688 2650 37088 6 Do0[1]
port 87 nsew signal output
rlabel metal2 s 53470 36688 53526 37088 6 Do0[20]
port 88 nsew signal output
rlabel metal2 s 55218 36688 55274 37088 6 Do0[21]
port 89 nsew signal output
rlabel metal2 s 56966 36688 57022 37088 6 Do0[22]
port 90 nsew signal output
rlabel metal2 s 58714 36688 58770 37088 6 Do0[23]
port 91 nsew signal output
rlabel metal2 s 60462 36688 60518 37088 6 Do0[24]
port 92 nsew signal output
rlabel metal2 s 62302 36688 62358 37088 6 Do0[25]
port 93 nsew signal output
rlabel metal2 s 64050 36688 64106 37088 6 Do0[26]
port 94 nsew signal output
rlabel metal2 s 65798 36688 65854 37088 6 Do0[27]
port 95 nsew signal output
rlabel metal2 s 67546 36688 67602 37088 6 Do0[28]
port 96 nsew signal output
rlabel metal2 s 69294 36688 69350 37088 6 Do0[29]
port 97 nsew signal output
rlabel metal2 s 4342 36688 4398 37088 6 Do0[2]
port 98 nsew signal output
rlabel metal2 s 71042 36688 71098 37088 6 Do0[30]
port 99 nsew signal output
rlabel metal2 s 72790 36688 72846 37088 6 Do0[31]
port 100 nsew signal output
rlabel metal2 s 74538 36688 74594 37088 6 Do0[32]
port 101 nsew signal output
rlabel metal2 s 76286 36688 76342 37088 6 Do0[33]
port 102 nsew signal output
rlabel metal2 s 78034 36688 78090 37088 6 Do0[34]
port 103 nsew signal output
rlabel metal2 s 79782 36688 79838 37088 6 Do0[35]
port 104 nsew signal output
rlabel metal2 s 81530 36688 81586 37088 6 Do0[36]
port 105 nsew signal output
rlabel metal2 s 83370 36688 83426 37088 6 Do0[37]
port 106 nsew signal output
rlabel metal2 s 85118 36688 85174 37088 6 Do0[38]
port 107 nsew signal output
rlabel metal2 s 86866 36688 86922 37088 6 Do0[39]
port 108 nsew signal output
rlabel metal2 s 6090 36688 6146 37088 6 Do0[3]
port 109 nsew signal output
rlabel metal2 s 88614 36688 88670 37088 6 Do0[40]
port 110 nsew signal output
rlabel metal2 s 90362 36688 90418 37088 6 Do0[41]
port 111 nsew signal output
rlabel metal2 s 92110 36688 92166 37088 6 Do0[42]
port 112 nsew signal output
rlabel metal2 s 93858 36688 93914 37088 6 Do0[43]
port 113 nsew signal output
rlabel metal2 s 95606 36688 95662 37088 6 Do0[44]
port 114 nsew signal output
rlabel metal2 s 97354 36688 97410 37088 6 Do0[45]
port 115 nsew signal output
rlabel metal2 s 99102 36688 99158 37088 6 Do0[46]
port 116 nsew signal output
rlabel metal2 s 100850 36688 100906 37088 6 Do0[47]
port 117 nsew signal output
rlabel metal2 s 102598 36688 102654 37088 6 Do0[48]
port 118 nsew signal output
rlabel metal2 s 104438 36688 104494 37088 6 Do0[49]
port 119 nsew signal output
rlabel metal2 s 7838 36688 7894 37088 6 Do0[4]
port 120 nsew signal output
rlabel metal2 s 106186 36688 106242 37088 6 Do0[50]
port 121 nsew signal output
rlabel metal2 s 107934 36688 107990 37088 6 Do0[51]
port 122 nsew signal output
rlabel metal2 s 109682 36688 109738 37088 6 Do0[52]
port 123 nsew signal output
rlabel metal2 s 111430 36688 111486 37088 6 Do0[53]
port 124 nsew signal output
rlabel metal2 s 113178 36688 113234 37088 6 Do0[54]
port 125 nsew signal output
rlabel metal2 s 114926 36688 114982 37088 6 Do0[55]
port 126 nsew signal output
rlabel metal2 s 116674 36688 116730 37088 6 Do0[56]
port 127 nsew signal output
rlabel metal2 s 118422 36688 118478 37088 6 Do0[57]
port 128 nsew signal output
rlabel metal2 s 120170 36688 120226 37088 6 Do0[58]
port 129 nsew signal output
rlabel metal2 s 121918 36688 121974 37088 6 Do0[59]
port 130 nsew signal output
rlabel metal2 s 9586 36688 9642 37088 6 Do0[5]
port 131 nsew signal output
rlabel metal2 s 123758 36688 123814 37088 6 Do0[60]
port 132 nsew signal output
rlabel metal2 s 125506 36688 125562 37088 6 Do0[61]
port 133 nsew signal output
rlabel metal2 s 127254 36688 127310 37088 6 Do0[62]
port 134 nsew signal output
rlabel metal2 s 129002 36688 129058 37088 6 Do0[63]
port 135 nsew signal output
rlabel metal2 s 11334 36688 11390 37088 6 Do0[6]
port 136 nsew signal output
rlabel metal2 s 13082 36688 13138 37088 6 Do0[7]
port 137 nsew signal output
rlabel metal2 s 14830 36688 14886 37088 6 Do0[8]
port 138 nsew signal output
rlabel metal2 s 16578 36688 16634 37088 6 Do0[9]
port 139 nsew signal output
rlabel metal2 s 20074 36688 20130 37088 6 Do1[0]
port 140 nsew signal output
rlabel metal2 s 130750 36688 130806 37088 6 Do1[10]
port 141 nsew signal output
rlabel metal2 s 132498 36688 132554 37088 6 Do1[11]
port 142 nsew signal output
rlabel metal2 s 134246 36688 134302 37088 6 Do1[12]
port 143 nsew signal output
rlabel metal2 s 135994 36688 136050 37088 6 Do1[13]
port 144 nsew signal output
rlabel metal2 s 137742 36688 137798 37088 6 Do1[14]
port 145 nsew signal output
rlabel metal2 s 139490 36688 139546 37088 6 Do1[15]
port 146 nsew signal output
rlabel metal2 s 141238 36688 141294 37088 6 Do1[16]
port 147 nsew signal output
rlabel metal2 s 142986 36688 143042 37088 6 Do1[17]
port 148 nsew signal output
rlabel metal2 s 144826 36688 144882 37088 6 Do1[18]
port 149 nsew signal output
rlabel metal2 s 146574 36688 146630 37088 6 Do1[19]
port 150 nsew signal output
rlabel metal2 s 23662 36688 23718 37088 6 Do1[1]
port 151 nsew signal output
rlabel metal2 s 148322 36688 148378 37088 6 Do1[20]
port 152 nsew signal output
rlabel metal2 s 150070 36688 150126 37088 6 Do1[21]
port 153 nsew signal output
rlabel metal2 s 151818 36688 151874 37088 6 Do1[22]
port 154 nsew signal output
rlabel metal2 s 153566 36688 153622 37088 6 Do1[23]
port 155 nsew signal output
rlabel metal2 s 155314 36688 155370 37088 6 Do1[24]
port 156 nsew signal output
rlabel metal2 s 157062 36688 157118 37088 6 Do1[25]
port 157 nsew signal output
rlabel metal2 s 158810 36688 158866 37088 6 Do1[26]
port 158 nsew signal output
rlabel metal2 s 160558 36688 160614 37088 6 Do1[27]
port 159 nsew signal output
rlabel metal2 s 162306 36688 162362 37088 6 Do1[28]
port 160 nsew signal output
rlabel metal2 s 164054 36688 164110 37088 6 Do1[29]
port 161 nsew signal output
rlabel metal2 s 27158 36688 27214 37088 6 Do1[2]
port 162 nsew signal output
rlabel metal2 s 165894 36688 165950 37088 6 Do1[30]
port 163 nsew signal output
rlabel metal2 s 167642 36688 167698 37088 6 Do1[31]
port 164 nsew signal output
rlabel metal2 s 169390 36688 169446 37088 6 Do1[32]
port 165 nsew signal output
rlabel metal2 s 171138 36688 171194 37088 6 Do1[33]
port 166 nsew signal output
rlabel metal2 s 172886 36688 172942 37088 6 Do1[34]
port 167 nsew signal output
rlabel metal2 s 174634 36688 174690 37088 6 Do1[35]
port 168 nsew signal output
rlabel metal2 s 176382 36688 176438 37088 6 Do1[36]
port 169 nsew signal output
rlabel metal2 s 178130 36688 178186 37088 6 Do1[37]
port 170 nsew signal output
rlabel metal2 s 179878 36688 179934 37088 6 Do1[38]
port 171 nsew signal output
rlabel metal2 s 181626 36688 181682 37088 6 Do1[39]
port 172 nsew signal output
rlabel metal2 s 30654 36688 30710 37088 6 Do1[3]
port 173 nsew signal output
rlabel metal2 s 183374 36688 183430 37088 6 Do1[40]
port 174 nsew signal output
rlabel metal2 s 185214 36688 185270 37088 6 Do1[41]
port 175 nsew signal output
rlabel metal2 s 186962 36688 187018 37088 6 Do1[42]
port 176 nsew signal output
rlabel metal2 s 188710 36688 188766 37088 6 Do1[43]
port 177 nsew signal output
rlabel metal2 s 190458 36688 190514 37088 6 Do1[44]
port 178 nsew signal output
rlabel metal2 s 192206 36688 192262 37088 6 Do1[45]
port 179 nsew signal output
rlabel metal2 s 193954 36688 194010 37088 6 Do1[46]
port 180 nsew signal output
rlabel metal2 s 195702 36688 195758 37088 6 Do1[47]
port 181 nsew signal output
rlabel metal2 s 197450 36688 197506 37088 6 Do1[48]
port 182 nsew signal output
rlabel metal2 s 199198 36688 199254 37088 6 Do1[49]
port 183 nsew signal output
rlabel metal2 s 34150 36688 34206 37088 6 Do1[4]
port 184 nsew signal output
rlabel metal2 s 200946 36688 201002 37088 6 Do1[50]
port 185 nsew signal output
rlabel metal2 s 202694 36688 202750 37088 6 Do1[51]
port 186 nsew signal output
rlabel metal2 s 204442 36688 204498 37088 6 Do1[52]
port 187 nsew signal output
rlabel metal2 s 206282 36688 206338 37088 6 Do1[53]
port 188 nsew signal output
rlabel metal2 s 208030 36688 208086 37088 6 Do1[54]
port 189 nsew signal output
rlabel metal2 s 209778 36688 209834 37088 6 Do1[55]
port 190 nsew signal output
rlabel metal2 s 211526 36688 211582 37088 6 Do1[56]
port 191 nsew signal output
rlabel metal2 s 213274 36688 213330 37088 6 Do1[57]
port 192 nsew signal output
rlabel metal2 s 215022 36688 215078 37088 6 Do1[58]
port 193 nsew signal output
rlabel metal2 s 216770 36688 216826 37088 6 Do1[59]
port 194 nsew signal output
rlabel metal2 s 37646 36688 37702 37088 6 Do1[5]
port 195 nsew signal output
rlabel metal2 s 218518 36688 218574 37088 6 Do1[60]
port 196 nsew signal output
rlabel metal2 s 220266 36688 220322 37088 6 Do1[61]
port 197 nsew signal output
rlabel metal2 s 222014 36688 222070 37088 6 Do1[62]
port 198 nsew signal output
rlabel metal2 s 223762 36688 223818 37088 6 Do1[63]
port 199 nsew signal output
rlabel metal2 s 41142 36688 41198 37088 6 Do1[6]
port 200 nsew signal output
rlabel metal2 s 44730 36688 44786 37088 6 Do1[7]
port 201 nsew signal output
rlabel metal2 s 48226 36688 48282 37088 6 Do1[8]
port 202 nsew signal output
rlabel metal2 s 51722 36688 51778 37088 6 Do1[9]
port 203 nsew signal output
rlabel metal3 s 224356 1232 224756 1352 6 EN0
port 204 nsew signal input
rlabel metal3 s 0 34416 400 34536 6 EN1
port 205 nsew signal input
rlabel metal4 s 19242 496 19862 36496 6 VGND
port 206 nsew ground input
rlabel metal4 s 55242 496 55862 36496 6 VGND
port 206 nsew ground input
rlabel metal4 s 91242 496 91862 36496 6 VGND
port 206 nsew ground input
rlabel metal4 s 127242 496 127862 36496 6 VGND
port 206 nsew ground input
rlabel metal4 s 163242 496 163862 36496 6 VGND
port 206 nsew ground input
rlabel metal4 s 199242 496 199862 36496 6 VGND
port 206 nsew ground input
rlabel metal4 s 1242 496 1862 36496 6 VPWR
port 207 nsew power input
rlabel metal4 s 37242 496 37862 36496 6 VPWR
port 207 nsew power input
rlabel metal4 s 73242 496 73862 36496 6 VPWR
port 207 nsew power input
rlabel metal4 s 109242 496 109862 36496 6 VPWR
port 207 nsew power input
rlabel metal4 s 145242 496 145862 36496 6 VPWR
port 207 nsew power input
rlabel metal4 s 181242 496 181862 36496 6 VPWR
port 207 nsew power input
rlabel metal4 s 217242 496 217862 36496 6 VPWR
port 207 nsew power input
rlabel metal3 s 224356 3816 224756 3936 6 WE0[0]
port 208 nsew signal input
rlabel metal3 s 224356 6536 224756 6656 6 WE0[1]
port 209 nsew signal input
rlabel metal3 s 224356 9120 224756 9240 6 WE0[2]
port 210 nsew signal input
rlabel metal3 s 224356 11840 224756 11960 6 WE0[3]
port 211 nsew signal input
rlabel metal3 s 224356 14424 224756 14544 6 WE0[4]
port 212 nsew signal input
rlabel metal3 s 224356 17144 224756 17264 6 WE0[5]
port 213 nsew signal input
rlabel metal3 s 224356 19728 224756 19848 6 WE0[6]
port 214 nsew signal input
rlabel metal3 s 224356 22448 224756 22568 6 WE0[7]
port 215 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 224756 37088
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17796730
string GDS_FILE /mnt/dffram/build/32x64_1RW1R/openlane/runs/RUN_2022.02.20_10.34.23/results/finishing/RAM32_1RW1R.magic.gds
string GDS_START 150134
<< end >>

