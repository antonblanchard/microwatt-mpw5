* NGSPICE file created from multiply_add_64x64.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_2 abstract view
.subckt sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_1 abstract view
.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_1 abstract view
.subckt sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_2 abstract view
.subckt sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_4 abstract view
.subckt sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

.subckt multiply_add_64x64 VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16]
+ a[17] a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29]
+ a[2] a[30] a[31] a[32] a[33] a[34] a[35] a[36] a[37] a[38] a[39] a[3] a[40] a[41]
+ a[42] a[43] a[44] a[45] a[46] a[47] a[48] a[49] a[4] a[50] a[51] a[52] a[53] a[54]
+ a[55] a[56] a[57] a[58] a[59] a[5] a[60] a[61] a[62] a[63] a[6] a[7] a[8] a[9] b[0]
+ b[10] b[11] b[12] b[13] b[14] b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22]
+ b[23] b[24] b[25] b[26] b[27] b[28] b[29] b[2] b[30] b[31] b[32] b[33] b[34] b[35]
+ b[36] b[37] b[38] b[39] b[3] b[40] b[41] b[42] b[43] b[44] b[45] b[46] b[47] b[48]
+ b[49] b[4] b[50] b[51] b[52] b[53] b[54] b[55] b[56] b[57] b[58] b[59] b[5] b[60]
+ b[61] b[62] b[63] b[6] b[7] b[8] b[9] c[0] c[100] c[101] c[102] c[103] c[104] c[105]
+ c[106] c[107] c[108] c[109] c[10] c[110] c[111] c[112] c[113] c[114] c[115] c[116]
+ c[117] c[118] c[119] c[11] c[120] c[121] c[122] c[123] c[124] c[125] c[126] c[127]
+ c[12] c[13] c[14] c[15] c[16] c[17] c[18] c[19] c[1] c[20] c[21] c[22] c[23] c[24]
+ c[25] c[26] c[27] c[28] c[29] c[2] c[30] c[31] c[32] c[33] c[34] c[35] c[36] c[37]
+ c[38] c[39] c[3] c[40] c[41] c[42] c[43] c[44] c[45] c[46] c[47] c[48] c[49] c[4]
+ c[50] c[51] c[52] c[53] c[54] c[55] c[56] c[57] c[58] c[59] c[5] c[60] c[61] c[62]
+ c[63] c[64] c[65] c[66] c[67] c[68] c[69] c[6] c[70] c[71] c[72] c[73] c[74] c[75]
+ c[76] c[77] c[78] c[79] c[7] c[80] c[81] c[82] c[83] c[84] c[85] c[86] c[87] c[88]
+ c[89] c[8] c[90] c[91] c[92] c[93] c[94] c[95] c[96] c[97] c[98] c[99] c[9] clk
+ o[0] o[100] o[101] o[102] o[103] o[104] o[105] o[106] o[107] o[108] o[109] o[10]
+ o[110] o[111] o[112] o[113] o[114] o[115] o[116] o[117] o[118] o[119] o[11] o[120]
+ o[121] o[122] o[123] o[124] o[125] o[126] o[127] o[12] o[13] o[14] o[15] o[16] o[17]
+ o[18] o[19] o[1] o[20] o[21] o[22] o[23] o[24] o[25] o[26] o[27] o[28] o[29] o[2]
+ o[30] o[31] o[32] o[33] o[34] o[35] o[36] o[37] o[38] o[39] o[3] o[40] o[41] o[42]
+ o[43] o[44] o[45] o[46] o[47] o[48] o[49] o[4] o[50] o[51] o[52] o[53] o[54] o[55]
+ o[56] o[57] o[58] o[59] o[5] o[60] o[61] o[62] o[63] o[64] o[65] o[66] o[67] o[68]
+ o[69] o[6] o[70] o[71] o[72] o[73] o[74] o[75] o[76] o[77] o[78] o[79] o[7] o[80]
+ o[81] o[82] o[83] o[84] o[85] o[86] o[87] o[88] o[89] o[8] o[90] o[91] o[92] o[93]
+ o[94] o[95] o[96] o[97] o[98] o[99] o[9] rst
XFILLER_140_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_57_8 dadda_fa_1_57_8/A dadda_fa_1_57_8/B dadda_fa_1_57_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_58_3/A dadda_fa_3_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_104_0 _695__915/HI U$$2875/X U$$3008/X VGND VGND VPWR VPWR dadda_fa_3_105_2/CIN
+ dadda_fa_3_104_3/B sky130_fd_sc_hd__fa_1
XFILLER_63_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1290 U$$1290/A U$$1342/B VGND VGND VPWR VPWR U$$1290/X sky130_fd_sc_hd__xor2_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_90_2 U$$2581/X U$$2714/X U$$2847/X VGND VGND VPWR VPWR dadda_fa_2_91_4/CIN
+ dadda_fa_2_90_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_1 U$$1769/X U$$1902/X U$$2035/X VGND VGND VPWR VPWR dadda_fa_2_84_2/A
+ dadda_fa_2_83_4/B sky130_fd_sc_hd__fa_2
XFILLER_172_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_60_0 dadda_fa_4_60_0/A dadda_fa_4_60_0/B dadda_fa_4_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/A dadda_fa_5_60_1/A sky130_fd_sc_hd__fa_1
XFILLER_172_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_76_0 U$$1489/X U$$1622/X U$$1755/X VGND VGND VPWR VPWR dadda_fa_2_77_0/B
+ dadda_fa_2_76_3/B sky130_fd_sc_hd__fa_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3609 U$$3609/A U$$3625/B VGND VGND VPWR VPWR U$$3609/X sky130_fd_sc_hd__xor2_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2908 U$$2908/A U$$2960/B VGND VGND VPWR VPWR U$$2908/X sky130_fd_sc_hd__xor2_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_501_ _501_/CLK _501_/D VGND VGND VPWR VPWR _501_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2919 U$$4289/A1 U$$2975/A2 U$$4289/B1 U$$2975/B2 VGND VGND VPWR VPWR U$$2920/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_5_124_1 U$$4511/X input156/X VGND VGND VPWR VPWR dadda_fa_6_125_0/CIN dadda_fa_7_124_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _432_/CLK _432_/D VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _632_/CLK _363_/D VGND VGND VPWR VPWR _363_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_294_ _612_/CLK _294_/D VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_98_1 dadda_fa_3_98_1/A dadda_fa_3_98_1/B dadda_fa_3_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_0/CIN dadda_fa_4_98_2/A sky130_fd_sc_hd__fa_1
XFILLER_5_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_75_0 dadda_fa_6_75_0/A dadda_fa_6_75_0/B dadda_fa_6_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_76_0/B dadda_fa_7_75_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$370 U$$94/B1 U$$278/X U$$96/B1 U$$279/X VGND VGND VPWR VPWR U$$371/A sky130_fd_sc_hd__a22o_1
XU$$381 U$$381/A _621_/Q VGND VGND VPWR VPWR U$$381/X sky130_fd_sc_hd__xor2_1
XU$$392 U$$940/A1 U$$278/X U$$942/A1 U$$279/X VGND VGND VPWR VPWR U$$393/A sky130_fd_sc_hd__a22o_1
XFILLER_178_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_0 U$$2853/X U$$2986/X U$$3119/X VGND VGND VPWR VPWR dadda_fa_3_94_0/B
+ dadda_fa_3_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_62_6 dadda_fa_1_62_6/A dadda_fa_1_62_6/B dadda_fa_1_62_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/B dadda_fa_2_62_5/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_55_5 U$$2777/X U$$2910/X U$$3043/X VGND VGND VPWR VPWR dadda_fa_2_56_2/A
+ dadda_fa_2_55_5/A sky130_fd_sc_hd__fa_1
XFILLER_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_48_4 U$$1699/X U$$1832/X U$$1965/X VGND VGND VPWR VPWR dadda_fa_2_49_2/B
+ dadda_fa_2_48_5/A sky130_fd_sc_hd__fa_1
XFILLER_43_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_2 dadda_fa_4_18_2/A dadda_fa_4_18_2/B dadda_ha_3_18_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_19_0/CIN dadda_fa_5_18_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_92_0 dadda_fa_7_92_0/A dadda_fa_7_92_0/B dadda_fa_7_92_0/CIN VGND VGND
+ VPWR VPWR _517_/D _388_/D sky130_fd_sc_hd__fa_1
XFILLER_155_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4107 U$$819/A1 U$$4107/A2 U$$4107/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4108/A
+ sky130_fd_sc_hd__a22o_1
XU$$4118 _552_/Q U$$4244/A2 U$$969/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4119/A sky130_fd_sc_hd__a22o_1
XU$$4129 U$$4129/A U$$4246/A VGND VGND VPWR VPWR U$$4129/X sky130_fd_sc_hd__xor2_1
XFILLER_59_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3406 U$$4502/A1 U$$3292/X U$$4504/A1 U$$3293/X VGND VGND VPWR VPWR U$$3407/A sky130_fd_sc_hd__a22o_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3417 U$$3417/A _665_/Q VGND VGND VPWR VPWR U$$3417/X sky130_fd_sc_hd__xor2_1
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3428 _667_/Q U$$3428/B VGND VGND VPWR VPWR U$$3428/X sky130_fd_sc_hd__and2_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3439 U$$14/A1 U$$3525/A2 _556_/Q U$$3525/B2 VGND VGND VPWR VPWR U$$3440/A sky130_fd_sc_hd__a22o_1
XFILLER_19_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2705 _599_/Q U$$2729/A2 U$$926/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2706/A sky130_fd_sc_hd__a22o_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2716 U$$2716/A _655_/Q VGND VGND VPWR VPWR U$$2716/X sky130_fd_sc_hd__xor2_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2727 U$$4508/A1 U$$2729/A2 U$$4510/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2728/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2738 U$$2738/A _655_/Q VGND VGND VPWR VPWR U$$2738/X sky130_fd_sc_hd__xor2_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2749 U$$2749/A U$$2797/B VGND VGND VPWR VPWR U$$2749/X sky130_fd_sc_hd__xor2_2
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_2 U$$845/X U$$978/X U$$1111/X VGND VGND VPWR VPWR dadda_fa_4_21_1/A
+ dadda_fa_4_20_2/B sky130_fd_sc_hd__fa_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _598_/CLK _415_/D VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_346_ _474_/CLK _346_/D VGND VGND VPWR VPWR _346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ _280_/CLK _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_72_5 dadda_fa_2_72_5/A dadda_fa_2_72_5/B dadda_fa_2_72_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_2/A dadda_fa_4_72_0/A sky130_fd_sc_hd__fa_2
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_65_4 dadda_fa_2_65_4/A dadda_fa_2_65_4/B dadda_fa_2_65_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/CIN dadda_fa_3_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_58_3 dadda_fa_2_58_3/A dadda_fa_2_58_3/B dadda_fa_2_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/B dadda_fa_3_58_3/B sky130_fd_sc_hd__fa_1
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3940 U$$787/B1 U$$3970/A2 U$$654/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3941/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_28_1 dadda_fa_5_28_1/A dadda_fa_5_28_1/B dadda_fa_5_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/B dadda_fa_7_28_0/A sky130_fd_sc_hd__fa_1
XU$$3951 U$$3951/A U$$3969/B VGND VGND VPWR VPWR U$$3951/X sky130_fd_sc_hd__xor2_1
XU$$3962 _611_/Q U$$3970/A2 U$$539/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3963/A sky130_fd_sc_hd__a22o_1
XU$$3973 _673_/Q VGND VGND VPWR VPWR U$$3973/Y sky130_fd_sc_hd__inv_1
XU$$3984 U$$3984/A U$$4044/B VGND VGND VPWR VPWR U$$3984/X sky130_fd_sc_hd__xor2_2
XU$$3995 _559_/Q U$$4045/A2 U$$4271/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$3996/A sky130_fd_sc_hd__a22o_1
XFILLER_52_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_102_1 dadda_fa_5_102_1/A dadda_fa_5_102_1/B dadda_fa_5_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/B dadda_fa_7_102_0/A sky130_fd_sc_hd__fa_2
XFILLER_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput264 _274_/Q VGND VGND VPWR VPWR o[106] sky130_fd_sc_hd__buf_2
Xoutput275 _284_/Q VGND VGND VPWR VPWR o[116] sky130_fd_sc_hd__buf_2
XFILLER_99_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput286 _294_/Q VGND VGND VPWR VPWR o[126] sky130_fd_sc_hd__buf_2
X_748__800 VGND VGND VPWR VPWR _748__800/HI U$$3294/A1 sky130_fd_sc_hd__conb_1
Xoutput297 _188_/Q VGND VGND VPWR VPWR o[20] sky130_fd_sc_hd__buf_2
XFILLER_102_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_60_3 U$$3186/X U$$3319/X U$$3452/X VGND VGND VPWR VPWR dadda_fa_2_61_1/B
+ dadda_fa_2_60_4/B sky130_fd_sc_hd__fa_1
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_53_2 U$$1177/X U$$1310/X U$$1443/X VGND VGND VPWR VPWR dadda_fa_2_54_1/A
+ dadda_fa_2_53_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_30_1 dadda_fa_4_30_1/A dadda_fa_4_30_1/B dadda_fa_4_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/B dadda_fa_5_30_1/B sky130_fd_sc_hd__fa_2
XFILLER_67_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_46_1 U$$498/X U$$631/X U$$764/X VGND VGND VPWR VPWR dadda_fa_2_47_2/A
+ dadda_fa_2_46_4/B sky130_fd_sc_hd__fa_2
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_23_0 dadda_fa_4_23_0/A dadda_fa_4_23_0/B dadda_fa_4_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/A dadda_fa_5_23_1/A sky130_fd_sc_hd__fa_1
XFILLER_82_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_39_0 U$$85/X U$$218/X U$$351/X VGND VGND VPWR VPWR dadda_fa_2_40_4/A dadda_fa_2_39_5/B
+ sky130_fd_sc_hd__fa_2
XFILLER_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_200_ _456_/CLK _200_/D VGND VGND VPWR VPWR _200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_75_3 dadda_fa_3_75_3/A dadda_fa_3_75_3/B dadda_fa_3_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/B dadda_fa_4_75_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_68_2 dadda_fa_3_68_2/A dadda_fa_3_68_2/B dadda_fa_3_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/A dadda_fa_4_68_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_38_0 dadda_fa_6_38_0/A dadda_fa_6_38_0/B dadda_fa_6_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_39_0/B dadda_fa_7_38_0/CIN sky130_fd_sc_hd__fa_1
XU$$3203 U$$50/B1 U$$3241/A2 U$$876/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3204/A sky130_fd_sc_hd__a22o_1
XU$$3214 U$$3214/A U$$3244/B VGND VGND VPWR VPWR U$$3214/X sky130_fd_sc_hd__xor2_1
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3225 U$$4045/B1 U$$3243/A2 U$$76/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3226/A sky130_fd_sc_hd__a22o_1
XU$$3236 U$$3236/A _663_/Q VGND VGND VPWR VPWR U$$3236/X sky130_fd_sc_hd__xor2_1
XU$$2502 U$$4283/A1 U$$2534/A2 U$$4285/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2503/A
+ sky130_fd_sc_hd__a22o_1
XU$$3247 _596_/Q U$$3155/X _597_/Q U$$3156/X VGND VGND VPWR VPWR U$$3248/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$18 _442_/Q _314_/Q VGND VGND VPWR VPWR final_adder.U$$513/B1 final_adder.U$$640/A
+ sky130_fd_sc_hd__ha_2
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$29 _453_/Q _325_/Q VGND VGND VPWR VPWR final_adder.U$$157/B1 final_adder.U$$651/A
+ sky130_fd_sc_hd__ha_1
XU$$2513 U$$2513/A U$$2533/B VGND VGND VPWR VPWR U$$2513/X sky130_fd_sc_hd__xor2_1
XU$$3258 U$$3258/A U$$3270/B VGND VGND VPWR VPWR U$$3258/X sky130_fd_sc_hd__xor2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2524 U$$880/A1 U$$2534/A2 _578_/Q U$$2534/B2 VGND VGND VPWR VPWR U$$2525/A sky130_fd_sc_hd__a22o_1
XU$$3269 _607_/Q U$$3155/X _608_/Q U$$3156/X VGND VGND VPWR VPWR U$$3270/A sky130_fd_sc_hd__a22o_1
XU$$2535 U$$2535/A U$$2585/B VGND VGND VPWR VPWR U$$2535/X sky130_fd_sc_hd__xor2_1
XU$$2546 _588_/Q U$$2584/A2 _589_/Q U$$2584/B2 VGND VGND VPWR VPWR U$$2547/A sky130_fd_sc_hd__a22o_1
XU$$1801 U$$979/A1 U$$1903/A2 U$$979/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1802/A sky130_fd_sc_hd__a22o_1
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2557 U$$2557/A U$$2603/A VGND VGND VPWR VPWR U$$2557/X sky130_fd_sc_hd__xor2_1
XFILLER_62_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1812 U$$1812/A U$$1918/A VGND VGND VPWR VPWR U$$1812/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2568 _599_/Q U$$2470/X _600_/Q U$$2471/X VGND VGND VPWR VPWR U$$2569/A sky130_fd_sc_hd__a22o_1
XU$$1823 U$$4289/A1 U$$1903/A2 U$$4289/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1824/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2579 U$$2579/A U$$2603/A VGND VGND VPWR VPWR U$$2579/X sky130_fd_sc_hd__xor2_1
XU$$1834 U$$1834/A U$$1872/B VGND VGND VPWR VPWR U$$1834/X sky130_fd_sc_hd__xor2_1
XU$$1845 U$$3900/A1 U$$1903/A2 U$$3489/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1846/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1856 U$$1856/A U$$1856/B VGND VGND VPWR VPWR U$$1856/X sky130_fd_sc_hd__xor2_1
XU$$1867 U$$771/A1 U$$1867/A2 U$$771/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1868/A sky130_fd_sc_hd__a22o_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1878 U$$1878/A U$$1904/B VGND VGND VPWR VPWR U$$1878/X sky130_fd_sc_hd__xor2_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1889 _602_/Q U$$1903/A2 _603_/Q U$$1903/B2 VGND VGND VPWR VPWR U$$1890/A sky130_fd_sc_hd__a22o_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_329_ _329_/CLK _329_/D VGND VGND VPWR VPWR _329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR _632_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_70_2 dadda_fa_2_70_2/A dadda_fa_2_70_2/B dadda_fa_2_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/A dadda_fa_3_70_3/A sky130_fd_sc_hd__fa_1
XFILLER_69_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_63_1 dadda_fa_2_63_1/A dadda_fa_2_63_1/B dadda_fa_2_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/CIN dadda_fa_3_63_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater701 U$$880/A1 VGND VGND VPWR VPWR U$$58/A1 sky130_fd_sc_hd__buf_12
XFILLER_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater712 _574_/Q VGND VGND VPWR VPWR U$$52/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$519 final_adder.U$$646/A final_adder.U$$646/B final_adder.U$$519/B1
+ VGND VGND VPWR VPWR final_adder.U$$647/B sky130_fd_sc_hd__a21o_1
XFILLER_56_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater723 _569_/Q VGND VGND VPWR VPWR U$$3876/B1 sky130_fd_sc_hd__buf_12
Xdadda_fa_5_40_0 dadda_fa_5_40_0/A dadda_fa_5_40_0/B dadda_fa_5_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/A dadda_fa_6_40_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_56_0 dadda_fa_2_56_0/A dadda_fa_2_56_0/B dadda_fa_2_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/B dadda_fa_3_56_2/B sky130_fd_sc_hd__fa_2
Xrepeater734 _564_/Q VGND VGND VPWR VPWR U$$32/A1 sky130_fd_sc_hd__buf_12
Xrepeater745 U$$842/A1 VGND VGND VPWR VPWR U$$20/A1 sky130_fd_sc_hd__buf_12
Xrepeater756 U$$4122/A1 VGND VGND VPWR VPWR U$$12/A1 sky130_fd_sc_hd__buf_12
XU$$4460 U$$759/B1 U$$4388/X U$$78/A1 U$$4389/X VGND VGND VPWR VPWR U$$4461/A sky130_fd_sc_hd__a22o_2
XU$$4471 U$$4471/A U$$4471/B VGND VGND VPWR VPWR U$$4471/X sky130_fd_sc_hd__xor2_1
XFILLER_93_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4482 U$$98/A1 U$$4388/X U$$4484/A1 U$$4389/X VGND VGND VPWR VPWR U$$4483/A sky130_fd_sc_hd__a22o_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4493 U$$4493/A U$$4493/B VGND VGND VPWR VPWR U$$4493/X sky130_fd_sc_hd__xor2_1
XFILLER_38_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3770 U$$3770/A U$$3794/B VGND VGND VPWR VPWR U$$3770/X sky130_fd_sc_hd__xor2_1
XU$$3781 U$$82/A1 U$$3783/A2 U$$632/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3782/A sky130_fd_sc_hd__a22o_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3792 U$$3792/A _671_/Q VGND VGND VPWR VPWR U$$3792/X sky130_fd_sc_hd__xor2_1
XFILLER_53_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_85_2 dadda_fa_4_85_2/A dadda_fa_4_85_2/B dadda_fa_4_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/CIN dadda_fa_5_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_78_1 dadda_fa_4_78_1/A dadda_fa_4_78_1/B dadda_fa_4_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/B dadda_fa_5_78_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_7_55_0 dadda_fa_7_55_0/A dadda_fa_7_55_0/B dadda_fa_7_55_0/CIN VGND VGND
+ VPWR VPWR _480_/D _351_/D sky130_fd_sc_hd__fa_1
XFILLER_121_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$903 U$$903/A U$$903/B VGND VGND VPWR VPWR U$$903/X sky130_fd_sc_hd__xor2_1
XU$$914 U$$914/A1 U$$928/A2 U$$92/B1 U$$928/B2 VGND VGND VPWR VPWR U$$915/A sky130_fd_sc_hd__a22o_1
XFILLER_29_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$925 U$$925/A U$$943/B VGND VGND VPWR VPWR U$$925/X sky130_fd_sc_hd__xor2_1
XFILLER_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$936 U$$936/A1 U$$826/X U$$938/A1 U$$827/X VGND VGND VPWR VPWR U$$937/A sky130_fd_sc_hd__a22o_1
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$947 U$$947/A _629_/Q VGND VGND VPWR VPWR U$$947/X sky130_fd_sc_hd__xor2_1
XU$$958 _629_/Q VGND VGND VPWR VPWR U$$958/Y sky130_fd_sc_hd__inv_1
XU$$969 U$$969/A1 U$$963/X U$$971/A1 U$$999/B2 VGND VGND VPWR VPWR U$$970/A sky130_fd_sc_hd__a22o_1
XU$$1108 U$$971/A1 U$$1100/X U$$12/B1 U$$1101/X VGND VGND VPWR VPWR U$$1109/A sky130_fd_sc_hd__a22o_1
XU$$1119 U$$1119/A U$$1189/B VGND VGND VPWR VPWR U$$1119/X sky130_fd_sc_hd__xor2_1
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_80_1 dadda_fa_3_80_1/A dadda_fa_3_80_1/B dadda_fa_3_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/CIN dadda_fa_4_80_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_0 dadda_fa_3_73_0/A dadda_fa_3_73_0/B dadda_fa_3_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/B dadda_fa_4_73_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_65_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3000 U$$3000/A U$$3004/B VGND VGND VPWR VPWR U$$3000/X sky130_fd_sc_hd__xor2_1
XFILLER_82_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3011 U$$956/A1 U$$2881/X U$$3011/B1 U$$2882/X VGND VGND VPWR VPWR U$$3012/A sky130_fd_sc_hd__a22o_1
XFILLER_93_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3022 U$$4255/A1 U$$3090/A2 _553_/Q U$$3090/B2 VGND VGND VPWR VPWR U$$3023/A sky130_fd_sc_hd__a22o_1
XFILLER_75_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3033 U$$3033/A U$$3085/B VGND VGND VPWR VPWR U$$3033/X sky130_fd_sc_hd__xor2_1
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3044 U$$30/A1 U$$3090/A2 U$$30/B1 U$$3090/B2 VGND VGND VPWR VPWR U$$3045/A sky130_fd_sc_hd__a22o_1
XU$$2310 U$$940/A1 U$$2316/A2 U$$942/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2311/A sky130_fd_sc_hd__a22o_1
XU$$3055 U$$3055/A U$$3085/B VGND VGND VPWR VPWR U$$3055/X sky130_fd_sc_hd__xor2_1
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_102_0 dadda_fa_4_102_0/A dadda_fa_4_102_0/B dadda_fa_4_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/A dadda_fa_5_102_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_35_5 U$$2338/X input185/X dadda_fa_2_35_5/CIN VGND VGND VPWR VPWR dadda_fa_3_36_2/A
+ dadda_fa_4_35_0/A sky130_fd_sc_hd__fa_2
XU$$3066 U$$52/A1 U$$3090/A2 U$$54/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3067/A sky130_fd_sc_hd__a22o_1
XU$$2321 U$$2321/A U$$2327/B VGND VGND VPWR VPWR U$$2321/X sky130_fd_sc_hd__xor2_1
XU$$3077 U$$3077/A U$$3137/B VGND VGND VPWR VPWR U$$3077/X sky130_fd_sc_hd__xor2_1
XU$$2332 U$$2464/B U$$2332/B VGND VGND VPWR VPWR U$$2332/X sky130_fd_sc_hd__and2_1
XFILLER_62_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2343 U$$12/B1 U$$2333/X U$$16/A1 U$$2334/X VGND VGND VPWR VPWR U$$2344/A sky130_fd_sc_hd__a22o_1
XU$$3088 _585_/Q U$$3018/X _586_/Q U$$3019/X VGND VGND VPWR VPWR U$$3089/A sky130_fd_sc_hd__a22o_1
XFILLER_61_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3099 U$$3099/A U$$3137/B VGND VGND VPWR VPWR U$$3099/X sky130_fd_sc_hd__xor2_1
XU$$2354 U$$2354/A U$$2432/B VGND VGND VPWR VPWR U$$2354/X sky130_fd_sc_hd__xor2_1
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1620 U$$1620/A U$$1643/A VGND VGND VPWR VPWR U$$1620/X sky130_fd_sc_hd__xor2_1
XU$$2365 U$$4283/A1 U$$2421/A2 U$$4285/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2366/A
+ sky130_fd_sc_hd__a22o_1
XU$$2376 U$$2376/A U$$2436/B VGND VGND VPWR VPWR U$$2376/X sky130_fd_sc_hd__xor2_1
XFILLER_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1631 _610_/Q U$$1641/A2 U$$4510/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1632/A sky130_fd_sc_hd__a22o_1
XU$$1642 U$$1642/A _639_/Q VGND VGND VPWR VPWR U$$1642/X sky130_fd_sc_hd__xor2_1
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2387 U$$880/A1 U$$2421/A2 _578_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2388/A sky130_fd_sc_hd__a22o_1
XU$$2398 U$$2398/A U$$2464/B VGND VGND VPWR VPWR U$$2398/X sky130_fd_sc_hd__xor2_1
XU$$1653 U$$1653/A U$$1781/A VGND VGND VPWR VPWR U$$1653/X sky130_fd_sc_hd__xor2_1
XU$$1664 U$$842/A1 U$$1734/A2 U$$22/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1665/A sky130_fd_sc_hd__a22o_1
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1675 U$$1675/A U$$1739/B VGND VGND VPWR VPWR U$$1675/X sky130_fd_sc_hd__xor2_1
XU$$1686 U$$3876/B1 U$$1726/A2 U$$4291/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1687/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1697 U$$1697/A U$$1727/B VGND VGND VPWR VPWR U$$1697/X sky130_fd_sc_hd__xor2_1
XFILLER_30_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_95_1 dadda_fa_5_95_1/A dadda_fa_5_95_1/B dadda_fa_5_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/B dadda_fa_7_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_88_0 dadda_fa_5_88_0/A dadda_fa_5_88_0/B dadda_fa_5_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/A dadda_fa_6_88_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_710__762 VGND VGND VPWR VPWR _710__762/HI U$$0/A sky130_fd_sc_hd__conb_1
XFILLER_85_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$305 final_adder.U$$304/A final_adder.U$$225/X final_adder.U$$227/X
+ VGND VGND VPWR VPWR final_adder.U$$305/X sky130_fd_sc_hd__a21o_1
XFILLER_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$316 final_adder.U$$316/A final_adder.U$$316/B VGND VGND VPWR VPWR
+ final_adder.U$$316/X sky130_fd_sc_hd__and2_1
XFILLER_85_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater520 _675_/Q VGND VGND VPWR VPWR U$$4044/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$327 final_adder.U$$326/A final_adder.U$$269/X final_adder.U$$271/X
+ VGND VGND VPWR VPWR final_adder.U$$327/X sky130_fd_sc_hd__a21o_1
Xrepeater531 _669_/Q VGND VGND VPWR VPWR U$$3625/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$338 final_adder.U$$338/A final_adder.U$$338/B VGND VGND VPWR VPWR
+ final_adder.U$$360/A sky130_fd_sc_hd__and2_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater542 U$$3129/B VGND VGND VPWR VPWR U$$3085/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$349 final_adder.U$$348/A final_adder.U$$313/X final_adder.U$$315/X
+ VGND VGND VPWR VPWR final_adder.U$$349/X sky130_fd_sc_hd__a21o_1
XFILLER_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater553 U$$2710/B VGND VGND VPWR VPWR U$$2698/B sky130_fd_sc_hd__buf_12
Xrepeater564 _647_/Q VGND VGND VPWR VPWR U$$2192/A sky130_fd_sc_hd__buf_12
Xrepeater575 U$$1739/B VGND VGND VPWR VPWR U$$1727/B sky130_fd_sc_hd__buf_12
Xrepeater586 _635_/Q VGND VGND VPWR VPWR U$$1369/A sky130_fd_sc_hd__buf_12
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater597 U$$822/A VGND VGND VPWR VPWR U$$784/B sky130_fd_sc_hd__buf_12
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4290 U$$4290/A U$$4332/B VGND VGND VPWR VPWR U$$4290/X sky130_fd_sc_hd__xor2_1
XFILLER_26_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_90_0 dadda_fa_4_90_0/A dadda_fa_4_90_0/B dadda_fa_4_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/A dadda_fa_5_90_1/A sky130_fd_sc_hd__fa_1
XFILLER_193_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_104_2 input134/X dadda_fa_3_104_2/B dadda_fa_3_104_2/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_105_1/A dadda_fa_4_104_2/B sky130_fd_sc_hd__fa_1
XFILLER_107_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_118_0 dadda_fa_6_118_0/A dadda_fa_6_118_0/B dadda_fa_6_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_119_0/B dadda_fa_7_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$700 U$$700/A U$$784/B VGND VGND VPWR VPWR U$$700/X sky130_fd_sc_hd__xor2_1
X_663_ _667_/CLK _663_/D VGND VGND VPWR VPWR _663_/Q sky130_fd_sc_hd__dfxtp_4
XU$$711 U$$26/A1 U$$689/X U$$987/A1 U$$817/B2 VGND VGND VPWR VPWR U$$712/A sky130_fd_sc_hd__a22o_1
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_38_3 dadda_fa_3_38_3/A dadda_fa_3_38_3/B dadda_fa_3_38_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/B dadda_fa_4_38_2/CIN sky130_fd_sc_hd__fa_2
XU$$722 U$$722/A U$$778/B VGND VGND VPWR VPWR U$$722/X sky130_fd_sc_hd__xor2_1
XU$$733 U$$48/A1 U$$817/A2 U$$50/A1 U$$785/B2 VGND VGND VPWR VPWR U$$734/A sky130_fd_sc_hd__a22o_1
XU$$744 U$$744/A U$$778/B VGND VGND VPWR VPWR U$$744/X sky130_fd_sc_hd__xor2_2
XU$$755 U$$70/A1 U$$817/A2 U$$70/B1 U$$785/B2 VGND VGND VPWR VPWR U$$756/A sky130_fd_sc_hd__a22o_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_594_ _594_/CLK _594_/D VGND VGND VPWR VPWR _594_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$766 U$$766/A U$$822/A VGND VGND VPWR VPWR U$$766/X sky130_fd_sc_hd__xor2_1
XU$$777 U$$92/A1 U$$785/A2 U$$92/B1 U$$785/B2 VGND VGND VPWR VPWR U$$778/A sky130_fd_sc_hd__a22o_1
XFILLER_72_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$788 U$$788/A U$$822/A VGND VGND VPWR VPWR U$$788/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$799 U$$799/A1 U$$689/X U$$938/A1 U$$690/X VGND VGND VPWR VPWR U$$800/A sky130_fd_sc_hd__a22o_1
XFILLER_188_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_700__920 VGND VGND VPWR VPWR _700__920/HI _700__920/LO sky130_fd_sc_hd__conb_1
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_40_3 U$$2747/X U$$2797/B input191/X VGND VGND VPWR VPWR dadda_fa_3_41_1/B
+ dadda_fa_3_40_3/B sky130_fd_sc_hd__fa_1
XFILLER_48_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_33_2 U$$871/X U$$1004/X U$$1137/X VGND VGND VPWR VPWR dadda_fa_3_34_1/A
+ dadda_fa_3_33_3/A sky130_fd_sc_hd__fa_1
X_699__919 VGND VGND VPWR VPWR _699__919/HI _699__919/LO sky130_fd_sc_hd__conb_1
XFILLER_23_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_10_1 dadda_fa_5_10_1/A dadda_fa_5_10_1/B dadda_ha_4_10_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_11_0/B dadda_fa_7_10_0/A sky130_fd_sc_hd__fa_2
XU$$2140 U$$2140/A _647_/Q VGND VGND VPWR VPWR U$$2140/X sky130_fd_sc_hd__xor2_1
XU$$2151 U$$96/A1 U$$2189/A2 U$$96/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2152/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_26_1 U$$458/X U$$591/X U$$724/X VGND VGND VPWR VPWR dadda_fa_3_27_2/CIN
+ dadda_fa_3_26_3/CIN sky130_fd_sc_hd__fa_2
XU$$2162 U$$2162/A U$$2192/A VGND VGND VPWR VPWR U$$2162/X sky130_fd_sc_hd__xor2_1
XFILLER_90_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2173 U$$940/A1 U$$2189/A2 U$$942/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2174/A sky130_fd_sc_hd__a22o_1
XU$$2184 U$$2184/A U$$2192/A VGND VGND VPWR VPWR U$$2184/X sky130_fd_sc_hd__xor2_1
XFILLER_62_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1450 U$$902/A1 U$$1472/A2 U$$902/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1451/A sky130_fd_sc_hd__a22o_1
XU$$2195 _649_/Q U$$2195/B VGND VGND VPWR VPWR U$$2195/X sky130_fd_sc_hd__and2_1
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1461 U$$1461/A U$$1461/B VGND VGND VPWR VPWR U$$1461/X sky130_fd_sc_hd__xor2_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1472 U$$924/A1 U$$1472/A2 U$$926/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1473/A sky130_fd_sc_hd__a22o_1
XU$$1483 U$$1483/A U$$1505/B VGND VGND VPWR VPWR U$$1483/X sky130_fd_sc_hd__xor2_1
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1494 U$$946/A1 U$$1374/X U$$948/A1 U$$1375/X VGND VGND VPWR VPWR U$$1495/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_85_5 U$$3502/X U$$3635/X U$$3768/X VGND VGND VPWR VPWR dadda_fa_2_86_4/A
+ dadda_fa_3_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_116_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_4 U$$2823/X U$$2956/X U$$3089/X VGND VGND VPWR VPWR dadda_fa_2_79_1/CIN
+ dadda_fa_2_78_4/CIN sky130_fd_sc_hd__fa_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$102 _526_/Q _398_/Q VGND VGND VPWR VPWR final_adder.U$$597/B1 final_adder.U$$724/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$113 _537_/Q _409_/Q VGND VGND VPWR VPWR final_adder.U$$241/B1 final_adder.U$$735/A
+ sky130_fd_sc_hd__ha_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$124 _548_/Q _420_/Q VGND VGND VPWR VPWR final_adder.U$$619/B1 final_adder.U$$746/A
+ sky130_fd_sc_hd__ha_1
XFILLER_44_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_48_2 dadda_fa_4_48_2/A dadda_fa_4_48_2/B dadda_fa_4_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/CIN dadda_fa_5_48_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$135 final_adder.U$$7/SUM final_adder.U$$6/COUT final_adder.U$$7/COUT
+ VGND VGND VPWR VPWR final_adder.U$$135/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$146 final_adder.U$$641/A final_adder.U$$640/A VGND VGND VPWR VPWR
+ final_adder.U$$264/A sky130_fd_sc_hd__and2_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$157 final_adder.U$$651/A final_adder.U$$523/B1 final_adder.U$$157/B1
+ VGND VGND VPWR VPWR final_adder.U$$157/X sky130_fd_sc_hd__a21o_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$168 final_adder.U$$663/A final_adder.U$$662/A VGND VGND VPWR VPWR
+ final_adder.U$$276/B sky130_fd_sc_hd__and2_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$179 final_adder.U$$673/A final_adder.U$$545/B1 final_adder.U$$179/B1
+ VGND VGND VPWR VPWR final_adder.U$$179/X sky130_fd_sc_hd__a21o_1
XFILLER_39_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater394 U$$4251/X VGND VGND VPWR VPWR U$$4381/A2 sky130_fd_sc_hd__buf_12
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_18_0 dadda_fa_7_18_0/A dadda_fa_7_18_0/B dadda_fa_7_18_0/CIN VGND VGND
+ VPWR VPWR _443_/D _314_/D sky130_fd_sc_hd__fa_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput120 b[5] VGND VGND VPWR VPWR _557_/D sky130_fd_sc_hd__clkbuf_4
Xinput131 c[101] VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__buf_4
Xdadda_fa_3_50_2 dadda_fa_3_50_2/A dadda_fa_3_50_2/B dadda_fa_3_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/A dadda_fa_4_50_2/B sky130_fd_sc_hd__fa_1
XFILLER_163_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput142 c[111] VGND VGND VPWR VPWR input142/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput153 c[121] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_0_66_2 U$$937/X U$$1070/X U$$1203/X VGND VGND VPWR VPWR dadda_fa_1_67_6/A
+ dadda_fa_1_66_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput164 c[16] VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput175 c[26] VGND VGND VPWR VPWR input175/X sky130_fd_sc_hd__buf_2
Xinput186 c[36] VGND VGND VPWR VPWR input186/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_43_1 dadda_fa_3_43_1/A dadda_fa_3_43_1/B dadda_fa_3_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/CIN dadda_fa_4_43_2/A sky130_fd_sc_hd__fa_2
Xdadda_fa_0_59_1 U$$524/X U$$657/X U$$790/X VGND VGND VPWR VPWR dadda_fa_1_60_6/CIN
+ dadda_fa_1_59_8/B sky130_fd_sc_hd__fa_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput197 c[46] VGND VGND VPWR VPWR input197/X sky130_fd_sc_hd__buf_4
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_20_0 dadda_fa_6_20_0/A dadda_fa_6_20_0/B dadda_fa_6_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_21_0/B dadda_fa_7_20_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$680 final_adder.U$$680/A final_adder.U$$680/B VGND VGND VPWR VPWR
+ _226_/D sky130_fd_sc_hd__xor2_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_36_0 dadda_fa_3_36_0/A dadda_fa_3_36_0/B dadda_fa_3_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/B dadda_fa_4_36_1/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$691 final_adder.U$$691/A final_adder.U$$691/B VGND VGND VPWR VPWR
+ _237_/D sky130_fd_sc_hd__xor2_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$530 U$$530/A U$$530/B VGND VGND VPWR VPWR U$$530/X sky130_fd_sc_hd__xor2_1
X_646_ _646_/CLK _646_/D VGND VGND VPWR VPWR _646_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$541 U$$952/A1 U$$415/X U$$952/B1 U$$416/X VGND VGND VPWR VPWR U$$542/A sky130_fd_sc_hd__a22o_1
XFILLER_17_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$552 U$$550/Y _624_/Q _623_/Q U$$551/X U$$548/Y VGND VGND VPWR VPWR U$$552/X sky130_fd_sc_hd__a32o_4
XFILLER_91_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$563 U$$563/A U$$661/B VGND VGND VPWR VPWR U$$563/X sky130_fd_sc_hd__xor2_1
XU$$574 U$$26/A1 U$$626/A2 U$$987/A1 U$$553/X VGND VGND VPWR VPWR U$$575/A sky130_fd_sc_hd__a22o_1
XFILLER_44_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$585 U$$585/A U$$623/B VGND VGND VPWR VPWR U$$585/X sky130_fd_sc_hd__xor2_1
XFILLER_60_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_577_ _578_/CLK _577_/D VGND VGND VPWR VPWR _577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$596 _572_/Q U$$626/A2 U$$735/A1 U$$553/X VGND VGND VPWR VPWR U$$597/A sky130_fd_sc_hd__a22o_1
XFILLER_108_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_95_4 U$$4187/X U$$4320/X U$$4453/X VGND VGND VPWR VPWR dadda_fa_3_96_1/CIN
+ dadda_fa_3_95_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_88_3 dadda_fa_2_88_3/A dadda_fa_2_88_3/B dadda_fa_2_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/B dadda_fa_3_88_3/B sky130_fd_sc_hd__fa_1
XFILLER_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_58_1 dadda_fa_5_58_1/A dadda_fa_5_58_1/B dadda_fa_5_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/B dadda_fa_7_58_0/A sky130_fd_sc_hd__fa_1
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_781__833 VGND VGND VPWR VPWR _781__833/HI U$$4407/B sky130_fd_sc_hd__conb_1
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_822__874 VGND VGND VPWR VPWR _822__874/HI U$$4489/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_104_1 U$$3141/X U$$3274/X U$$3407/X VGND VGND VPWR VPWR dadda_fa_3_105_3/A
+ dadda_fa_3_104_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1280 U$$1280/A U$$1342/B VGND VGND VPWR VPWR U$$1280/X sky130_fd_sc_hd__xor2_1
XU$$1291 U$$880/A1 U$$1341/A2 U$$4170/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1292/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_125_0 U$$4246/Y U$$4380/X U$$4513/X VGND VGND VPWR VPWR dadda_fa_6_126_0/CIN
+ dadda_fa_7_125_0/A sky130_fd_sc_hd__fa_2
XFILLER_164_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_2 U$$2168/X U$$2301/X U$$2434/X VGND VGND VPWR VPWR dadda_fa_2_84_2/B
+ dadda_fa_2_83_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_46_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_60_1 dadda_fa_4_60_1/A dadda_fa_4_60_1/B dadda_fa_4_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/B dadda_fa_5_60_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_76_1 U$$1888/X U$$2021/X U$$2154/X VGND VGND VPWR VPWR dadda_fa_2_77_0/CIN
+ dadda_fa_2_76_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_120_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_53_0 dadda_fa_4_53_0/A dadda_fa_4_53_0/B dadda_fa_4_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/A dadda_fa_5_53_1/A sky130_fd_sc_hd__fa_1
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_69_0 U$$2406/X U$$2539/X U$$2672/X VGND VGND VPWR VPWR dadda_fa_2_70_0/B
+ dadda_fa_2_69_3/B sky130_fd_sc_hd__fa_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_500_ _500_/CLK _500_/D VGND VGND VPWR VPWR _500_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2909 U$$32/A1 U$$3009/A2 U$$34/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2910/A sky130_fd_sc_hd__a22o_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_431_ _431_/CLK _431_/D VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _367_/CLK _362_/D VGND VGND VPWR VPWR _362_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_293_ _612_/CLK _293_/D VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_98_2 dadda_fa_3_98_2/A dadda_fa_3_98_2/B dadda_fa_3_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/A dadda_fa_4_98_2/B sky130_fd_sc_hd__fa_2
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_68_0 dadda_fa_6_68_0/A dadda_fa_6_68_0/B dadda_fa_6_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_69_0/B dadda_fa_7_68_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_765__817 VGND VGND VPWR VPWR _765__817/HI U$$4253/A1 sky130_fd_sc_hd__conb_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_71_0 U$$547/Y U$$681/X U$$814/X VGND VGND VPWR VPWR dadda_fa_1_72_6/CIN
+ dadda_fa_1_71_8/A sky130_fd_sc_hd__fa_1
XFILLER_7_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_806__858 VGND VGND VPWR VPWR _806__858/HI U$$4457/B sky130_fd_sc_hd__conb_1
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_5_7_1 U$$420/X input234/X VGND VGND VPWR VPWR dadda_fa_6_8_0/B dadda_fa_7_7_0/A
+ sky130_fd_sc_hd__ha_2
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$360 U$$86/A1 U$$278/X U$$88/A1 U$$279/X VGND VGND VPWR VPWR U$$361/A sky130_fd_sc_hd__a22o_1
X_629_ _633_/CLK _629_/D VGND VGND VPWR VPWR _629_/Q sky130_fd_sc_hd__dfxtp_4
XU$$371 U$$371/A U$$391/B VGND VGND VPWR VPWR U$$371/X sky130_fd_sc_hd__xor2_1
XFILLER_17_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$382 U$$930/A1 U$$278/X U$$932/A1 U$$279/X VGND VGND VPWR VPWR U$$383/A sky130_fd_sc_hd__a22o_1
XU$$393 U$$393/A _621_/Q VGND VGND VPWR VPWR U$$393/X sky130_fd_sc_hd__xor2_1
XFILLER_177_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_93_1 U$$3252/X U$$3385/X U$$3518/X VGND VGND VPWR VPWR dadda_fa_3_94_0/CIN
+ dadda_fa_3_93_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_70_0 dadda_fa_5_70_0/A dadda_fa_5_70_0/B dadda_fa_5_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/A dadda_fa_6_70_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_86_0 U$$3770/X U$$3903/X U$$4036/X VGND VGND VPWR VPWR dadda_fa_3_87_0/B
+ dadda_fa_3_86_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_1_49_7 U$$2898/X U$$3031/X VGND VGND VPWR VPWR dadda_fa_2_50_3/A dadda_fa_3_49_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_62_7 dadda_fa_1_62_7/A dadda_fa_1_62_7/B dadda_fa_1_62_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/CIN dadda_fa_2_62_5/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_1_55_6 U$$3176/X U$$3309/X U$$3442/X VGND VGND VPWR VPWR dadda_fa_2_56_2/B
+ dadda_fa_2_55_5/B sky130_fd_sc_hd__fa_1
XFILLER_83_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_48_5 U$$2098/X U$$2231/X U$$2364/X VGND VGND VPWR VPWR dadda_fa_2_49_2/CIN
+ dadda_fa_2_48_5/B sky130_fd_sc_hd__fa_1
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_7_0 dadda_fa_7_7_0/A dadda_fa_7_7_0/B dadda_fa_7_7_0/CIN VGND VGND VPWR
+ VPWR _432_/D _303_/D sky130_fd_sc_hd__fa_1
XFILLER_169_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_85_0 dadda_fa_7_85_0/A dadda_fa_7_85_0/B dadda_fa_7_85_0/CIN VGND VGND
+ VPWR VPWR _510_/D _381_/D sky130_fd_sc_hd__fa_2
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4108 U$$4108/A U$$4109/A VGND VGND VPWR VPWR U$$4108/X sky130_fd_sc_hd__xor2_1
XU$$4119 U$$4119/A _677_/Q VGND VGND VPWR VPWR U$$4119/X sky130_fd_sc_hd__xor2_1
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3407 U$$3407/A _665_/Q VGND VGND VPWR VPWR U$$3407/X sky130_fd_sc_hd__xor2_1
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3418 U$$4514/A1 U$$3292/X U$$4379/A1 U$$3293/X VGND VGND VPWR VPWR U$$3419/A sky130_fd_sc_hd__a22o_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3429 U$$3427/Y _666_/Q _665_/Q U$$3428/X U$$3425/Y VGND VGND VPWR VPWR U$$3429/X
+ sky130_fd_sc_hd__a32o_4
Xdadda_fa_6_100_0 dadda_fa_6_100_0/A dadda_fa_6_100_0/B dadda_fa_6_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_101_0/B dadda_fa_7_100_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2706 U$$2706/A U$$2710/B VGND VGND VPWR VPWR U$$2706/X sky130_fd_sc_hd__xor2_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2717 _605_/Q U$$2607/X _606_/Q U$$2608/X VGND VGND VPWR VPWR U$$2718/A sky130_fd_sc_hd__a22o_1
XFILLER_34_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2728 U$$2728/A _655_/Q VGND VGND VPWR VPWR U$$2728/X sky130_fd_sc_hd__xor2_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2739 _655_/Q VGND VGND VPWR VPWR U$$2739/Y sky130_fd_sc_hd__inv_1
XFILLER_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _594_/CLK _414_/D VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _483_/CLK _345_/D VGND VGND VPWR VPWR _345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_276_ _280_/CLK _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_65_5 dadda_fa_2_65_5/A dadda_fa_2_65_5/B dadda_fa_2_65_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_2/A dadda_fa_4_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_1_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_58_4 dadda_fa_2_58_4/A dadda_fa_2_58_4/B dadda_fa_2_58_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/CIN dadda_fa_3_58_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3930 U$$94/A1 U$$3970/A2 _596_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3931/A sky130_fd_sc_hd__a22o_1
XU$$3941 U$$3941/A _673_/Q VGND VGND VPWR VPWR U$$3941/X sky130_fd_sc_hd__xor2_1
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3952 U$$4500/A1 U$$3970/A2 U$$4502/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3953/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3963 U$$3963/A _673_/Q VGND VGND VPWR VPWR U$$3963/X sky130_fd_sc_hd__xor2_1
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3974 _674_/Q VGND VGND VPWR VPWR U$$3976/B sky130_fd_sc_hd__inv_1
XFILLER_18_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3985 U$$12/A1 U$$4045/A2 _555_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$3986/A sky130_fd_sc_hd__a22o_1
XFILLER_75_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3996 U$$3996/A U$$4044/B VGND VGND VPWR VPWR U$$3996/X sky130_fd_sc_hd__xor2_1
XFILLER_80_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$190 U$$190/A U$$262/B VGND VGND VPWR VPWR U$$190/X sky130_fd_sc_hd__xor2_1
XFILLER_178_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput265 _275_/Q VGND VGND VPWR VPWR o[107] sky130_fd_sc_hd__buf_2
XFILLER_160_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput276 _285_/Q VGND VGND VPWR VPWR o[117] sky130_fd_sc_hd__buf_2
XFILLER_0_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput287 _295_/Q VGND VGND VPWR VPWR o[127] sky130_fd_sc_hd__buf_2
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput298 _189_/Q VGND VGND VPWR VPWR o[21] sky130_fd_sc_hd__buf_2
XFILLER_102_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_60_4 U$$3585/X U$$3718/X U$$3851/X VGND VGND VPWR VPWR dadda_fa_2_61_1/CIN
+ dadda_fa_2_60_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_828__880 VGND VGND VPWR VPWR _828__880/HI U$$4501/B sky130_fd_sc_hd__conb_1
XFILLER_56_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_53_3 U$$1576/X U$$1709/X U$$1842/X VGND VGND VPWR VPWR dadda_fa_2_54_1/B
+ dadda_fa_2_53_4/B sky130_fd_sc_hd__fa_1
XFILLER_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_94_clk _632_/CLK VGND VGND VPWR VPWR _622_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_4_30_2 dadda_fa_4_30_2/A dadda_fa_4_30_2/B dadda_fa_4_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/CIN dadda_fa_5_30_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_46_2 U$$897/X U$$1030/X U$$1163/X VGND VGND VPWR VPWR dadda_fa_2_47_2/B
+ dadda_fa_2_46_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_167_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_23_1 dadda_fa_4_23_1/A dadda_fa_4_23_1/B dadda_fa_4_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/B dadda_fa_5_23_1/B sky130_fd_sc_hd__fa_2
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_39_1 U$$484/X U$$617/X U$$750/X VGND VGND VPWR VPWR dadda_fa_2_40_4/B
+ dadda_fa_2_39_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_16_0 U$$704/X U$$837/X U$$970/X VGND VGND VPWR VPWR dadda_fa_5_17_0/A
+ dadda_fa_5_16_1/A sky130_fd_sc_hd__fa_2
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_68_3 dadda_fa_3_68_3/A dadda_fa_3_68_3/B dadda_fa_3_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/B dadda_fa_4_68_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3204 U$$3204/A U$$3224/B VGND VGND VPWR VPWR U$$3204/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3215 U$$3900/A1 U$$3241/A2 U$$3489/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3216/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_85_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _642_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3226 U$$3226/A U$$3244/B VGND VGND VPWR VPWR U$$3226/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$19 _443_/Q _315_/Q VGND VGND VPWR VPWR final_adder.U$$147/B1 final_adder.U$$641/A
+ sky130_fd_sc_hd__ha_1
XU$$3237 U$$771/A1 U$$3241/A2 U$$771/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3238/A sky130_fd_sc_hd__a22o_1
XU$$2503 U$$2503/A U$$2533/B VGND VGND VPWR VPWR U$$2503/X sky130_fd_sc_hd__xor2_1
XU$$3248 U$$3248/A U$$3270/B VGND VGND VPWR VPWR U$$3248/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2514 U$$4156/B1 U$$2584/A2 _573_/Q U$$2584/B2 VGND VGND VPWR VPWR U$$2515/A sky130_fd_sc_hd__a22o_1
XFILLER_74_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3259 U$$928/B1 U$$3155/X U$$4494/A1 U$$3156/X VGND VGND VPWR VPWR U$$3260/A sky130_fd_sc_hd__a22o_1
XU$$2525 U$$2525/A U$$2585/B VGND VGND VPWR VPWR U$$2525/X sky130_fd_sc_hd__xor2_1
XFILLER_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2536 U$$892/A1 U$$2584/A2 U$$892/B1 U$$2584/B2 VGND VGND VPWR VPWR U$$2537/A sky130_fd_sc_hd__a22o_1
XU$$2547 U$$2547/A U$$2585/B VGND VGND VPWR VPWR U$$2547/X sky130_fd_sc_hd__xor2_1
XU$$1802 U$$1802/A U$$1856/B VGND VGND VPWR VPWR U$$1802/X sky130_fd_sc_hd__xor2_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1813 U$$30/B1 U$$1867/A2 U$$3457/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1814/A sky130_fd_sc_hd__a22o_1
XFILLER_27_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2558 U$$92/A1 U$$2584/A2 U$$92/B1 U$$2584/B2 VGND VGND VPWR VPWR U$$2559/A sky130_fd_sc_hd__a22o_1
XU$$2569 U$$2569/A U$$2603/A VGND VGND VPWR VPWR U$$2569/X sky130_fd_sc_hd__xor2_1
XU$$1824 U$$1824/A U$$1856/B VGND VGND VPWR VPWR U$$1824/X sky130_fd_sc_hd__xor2_1
XFILLER_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1835 U$$54/A1 U$$1867/A2 U$$56/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1836/A sky130_fd_sc_hd__a22o_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1846 U$$1846/A U$$1856/B VGND VGND VPWR VPWR U$$1846/X sky130_fd_sc_hd__xor2_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1857 U$$759/B1 U$$1867/A2 U$$78/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1858/A sky130_fd_sc_hd__a22o_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1868 U$$1868/A U$$1918/A VGND VGND VPWR VPWR U$$1868/X sky130_fd_sc_hd__xor2_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1879 _597_/Q U$$1903/A2 _598_/Q U$$1903/B2 VGND VGND VPWR VPWR U$$1880/A sky130_fd_sc_hd__a22o_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_328_ _329_/CLK _328_/D VGND VGND VPWR VPWR _328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_259_ _267_/CLK _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_3 dadda_fa_2_70_3/A dadda_fa_2_70_3/B dadda_fa_2_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/B dadda_fa_3_70_3/B sky130_fd_sc_hd__fa_1
XFILLER_124_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_63_2 dadda_fa_2_63_2/A dadda_fa_2_63_2/B dadda_fa_2_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/A dadda_fa_3_63_3/A sky130_fd_sc_hd__fa_2
XFILLER_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater702 U$$4442/A1 VGND VGND VPWR VPWR U$$880/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$509 final_adder.U$$636/A final_adder.U$$636/B final_adder.U$$509/B1
+ VGND VGND VPWR VPWR final_adder.U$$637/B sky130_fd_sc_hd__a21o_1
Xrepeater713 _573_/Q VGND VGND VPWR VPWR U$$50/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_5_40_1 dadda_fa_5_40_1/A dadda_fa_5_40_1/B dadda_fa_5_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/B dadda_fa_7_40_0/A sky130_fd_sc_hd__fa_2
Xrepeater724 U$$4424/A1 VGND VGND VPWR VPWR U$$3191/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_56_1 dadda_fa_2_56_1/A dadda_fa_2_56_1/B dadda_fa_2_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/CIN dadda_fa_3_56_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater735 U$$30/A1 VGND VGND VPWR VPWR U$$28/B1 sky130_fd_sc_hd__buf_12
XFILLER_84_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater746 U$$842/A1 VGND VGND VPWR VPWR U$$979/A1 sky130_fd_sc_hd__buf_12
XFILLER_42_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_33_0 dadda_fa_5_33_0/A dadda_fa_5_33_0/B dadda_fa_5_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/A dadda_fa_6_33_0/CIN sky130_fd_sc_hd__fa_2
Xrepeater757 _554_/Q VGND VGND VPWR VPWR U$$4122/A1 sky130_fd_sc_hd__buf_12
XU$$4450 _581_/Q U$$4388/X _582_/Q U$$4389/X VGND VGND VPWR VPWR U$$4451/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_76_clk _560_/CLK VGND VGND VPWR VPWR _656_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4461 U$$4461/A U$$4461/B VGND VGND VPWR VPWR U$$4461/X sky130_fd_sc_hd__xor2_4
Xdadda_fa_2_49_0 U$$3164/X U$$3297/X input200/X VGND VGND VPWR VPWR dadda_fa_3_50_0/B
+ dadda_fa_3_49_2/B sky130_fd_sc_hd__fa_2
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4472 U$$771/B1 U$$4388/X U$$90/A1 U$$4389/X VGND VGND VPWR VPWR U$$4473/A sky130_fd_sc_hd__a22o_2
XU$$4483 U$$4483/A U$$4483/B VGND VGND VPWR VPWR U$$4483/X sky130_fd_sc_hd__xor2_1
XU$$4494 U$$4494/A1 U$$4388/X U$$4496/A1 U$$4389/X VGND VGND VPWR VPWR U$$4495/A sky130_fd_sc_hd__a22o_1
XU$$3760 U$$3760/A U$$3784/B VGND VGND VPWR VPWR U$$3760/X sky130_fd_sc_hd__xor2_1
XU$$3771 U$$72/A1 U$$3795/A2 U$$4045/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3772/A sky130_fd_sc_hd__a22o_1
XU$$3782 U$$3782/A U$$3784/B VGND VGND VPWR VPWR U$$3782/X sky130_fd_sc_hd__xor2_1
XU$$3793 U$$94/A1 U$$3703/X _596_/Q U$$3704/X VGND VGND VPWR VPWR U$$3794/A sky130_fd_sc_hd__a22o_1
XFILLER_178_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_78_2 dadda_fa_4_78_2/A dadda_fa_4_78_2/B dadda_fa_4_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/CIN dadda_fa_5_78_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_48_0 dadda_fa_7_48_0/A dadda_fa_7_48_0/B dadda_fa_7_48_0/CIN VGND VGND
+ VPWR VPWR _473_/D _344_/D sky130_fd_sc_hd__fa_2
XFILLER_85_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_51_0 U$$109/X U$$242/X U$$375/X VGND VGND VPWR VPWR dadda_fa_2_52_0/B
+ dadda_fa_2_51_3/B sky130_fd_sc_hd__fa_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _581_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$904 U$$82/A1 U$$910/A2 U$$84/A1 U$$910/B2 VGND VGND VPWR VPWR U$$905/A sky130_fd_sc_hd__a22o_1
XFILLER_56_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$915 U$$915/A U$$943/B VGND VGND VPWR VPWR U$$915/X sky130_fd_sc_hd__xor2_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$926 U$$926/A1 U$$928/A2 U$$928/A1 U$$928/B2 VGND VGND VPWR VPWR U$$927/A sky130_fd_sc_hd__a22o_1
XU$$937 U$$937/A U$$943/B VGND VGND VPWR VPWR U$$937/X sky130_fd_sc_hd__xor2_1
XFILLER_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$948 U$$948/A1 U$$826/X U$$950/A1 U$$827/X VGND VGND VPWR VPWR U$$949/A sky130_fd_sc_hd__a22o_1
XU$$959 U$$959/A VGND VGND VPWR VPWR U$$959/Y sky130_fd_sc_hd__inv_1
XFILLER_16_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1109 U$$1109/A U$$1189/B VGND VGND VPWR VPWR U$$1109/X sky130_fd_sc_hd__xor2_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_2 dadda_fa_3_80_2/A dadda_fa_3_80_2/B dadda_fa_3_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/A dadda_fa_4_80_2/B sky130_fd_sc_hd__fa_2
XFILLER_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_73_1 dadda_fa_3_73_1/A dadda_fa_3_73_1/B dadda_fa_3_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/CIN dadda_fa_4_73_2/A sky130_fd_sc_hd__fa_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_50_0 dadda_fa_6_50_0/A dadda_fa_6_50_0/B dadda_fa_6_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_51_0/B dadda_fa_7_50_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_66_0 dadda_fa_3_66_0/A dadda_fa_3_66_0/B dadda_fa_3_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/B dadda_fa_4_66_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_182_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3001 U$$4508/A1 U$$2881/X _611_/Q U$$2882/X VGND VGND VPWR VPWR U$$3002/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_58_clk _536_/CLK VGND VGND VPWR VPWR _531_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3012 U$$3012/A _659_/Q VGND VGND VPWR VPWR U$$3012/X sky130_fd_sc_hd__xor2_1
XU$$3023 U$$3023/A U$$3085/B VGND VGND VPWR VPWR U$$3023/X sky130_fd_sc_hd__xor2_1
XU$$3034 U$$979/A1 U$$3090/A2 U$$979/B1 U$$3090/B2 VGND VGND VPWR VPWR U$$3035/A sky130_fd_sc_hd__a22o_1
XFILLER_75_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2300 _602_/Q U$$2326/A2 _603_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2301/A sky130_fd_sc_hd__a22o_1
XU$$3045 U$$3045/A U$$3085/B VGND VGND VPWR VPWR U$$3045/X sky130_fd_sc_hd__xor2_1
XU$$2311 U$$2311/A _649_/Q VGND VGND VPWR VPWR U$$2311/X sky130_fd_sc_hd__xor2_1
XU$$3056 U$$3876/B1 U$$3090/A2 U$$4291/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3057/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_102_1 dadda_fa_4_102_1/A dadda_fa_4_102_1/B dadda_fa_4_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/B dadda_fa_5_102_1/B sky130_fd_sc_hd__fa_1
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2322 U$$4514/A1 U$$2326/A2 U$$4379/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2323/A
+ sky130_fd_sc_hd__a22o_1
XU$$3067 U$$3067/A U$$3129/B VGND VGND VPWR VPWR U$$3067/X sky130_fd_sc_hd__xor2_1
XU$$3078 _580_/Q U$$3018/X _581_/Q U$$3019/X VGND VGND VPWR VPWR U$$3079/A sky130_fd_sc_hd__a22o_1
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2333 U$$2331/Y _650_/Q _649_/Q U$$2332/X U$$2329/Y VGND VGND VPWR VPWR U$$2333/X
+ sky130_fd_sc_hd__a32o_4
XU$$3089 U$$3089/A U$$3137/B VGND VGND VPWR VPWR U$$3089/X sky130_fd_sc_hd__xor2_1
XU$$2344 U$$2344/A U$$2432/B VGND VGND VPWR VPWR U$$2344/X sky130_fd_sc_hd__xor2_1
XU$$2355 U$$4273/A1 U$$2421/A2 U$$28/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2356/A sky130_fd_sc_hd__a22o_1
XFILLER_35_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1610 U$$1610/A U$$1614/B VGND VGND VPWR VPWR U$$1610/X sky130_fd_sc_hd__xor2_1
XFILLER_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1621 U$$936/A1 U$$1641/A2 _606_/Q U$$1641/B2 VGND VGND VPWR VPWR U$$1622/A sky130_fd_sc_hd__a22o_1
XU$$2366 U$$2366/A U$$2432/B VGND VGND VPWR VPWR U$$2366/X sky130_fd_sc_hd__xor2_1
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1632 U$$1632/A U$$1643/A VGND VGND VPWR VPWR U$$1632/X sky130_fd_sc_hd__xor2_1
XU$$2377 U$$48/A1 U$$2421/A2 U$$50/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2378/A sky130_fd_sc_hd__a22o_1
XU$$1643 U$$1643/A VGND VGND VPWR VPWR U$$1643/Y sky130_fd_sc_hd__inv_1
XU$$2388 U$$2388/A U$$2432/B VGND VGND VPWR VPWR U$$2388/X sky130_fd_sc_hd__xor2_1
XFILLER_188_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2399 U$$70/A1 U$$2333/X U$$70/B1 U$$2334/X VGND VGND VPWR VPWR U$$2400/A sky130_fd_sc_hd__a22o_1
XU$$1654 U$$8/B1 U$$1734/A2 U$$12/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1655/A sky130_fd_sc_hd__a22o_1
XU$$1665 U$$1665/A U$$1781/A VGND VGND VPWR VPWR U$$1665/X sky130_fd_sc_hd__xor2_1
XU$$1676 U$$32/A1 U$$1734/A2 U$$34/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1677/A sky130_fd_sc_hd__a22o_1
XFILLER_43_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1687 U$$1687/A U$$1727/B VGND VGND VPWR VPWR U$$1687/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_123_0 dadda_fa_7_123_0/A dadda_fa_7_123_0/B dadda_fa_7_123_0/CIN VGND
+ VGND VPWR VPWR _548_/D _419_/D sky130_fd_sc_hd__fa_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1698 U$$876/A1 U$$1726/A2 U$$878/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1699/A sky130_fd_sc_hd__a22o_1
XFILLER_148_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_88_1 dadda_fa_5_88_1/A dadda_fa_5_88_1/B dadda_fa_5_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/B dadda_fa_7_88_0/A sky130_fd_sc_hd__fa_2
XFILLER_115_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$306 final_adder.U$$306/A final_adder.U$$306/B VGND VGND VPWR VPWR
+ final_adder.U$$344/A sky130_fd_sc_hd__and2_1
Xrepeater510 U$$1375/X VGND VGND VPWR VPWR U$$1466/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$317 final_adder.U$$316/A final_adder.U$$249/X final_adder.U$$251/X
+ VGND VGND VPWR VPWR final_adder.U$$317/X sky130_fd_sc_hd__a21o_1
Xrepeater521 _675_/Q VGND VGND VPWR VPWR U$$4109/A sky130_fd_sc_hd__buf_12
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$328 final_adder.U$$328/A final_adder.U$$328/B VGND VGND VPWR VPWR
+ final_adder.U$$356/B sky130_fd_sc_hd__and2_1
Xrepeater532 _669_/Q VGND VGND VPWR VPWR U$$3699/A sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$339 final_adder.U$$338/A final_adder.U$$293/X final_adder.U$$295/X
+ VGND VGND VPWR VPWR final_adder.U$$339/X sky130_fd_sc_hd__a21o_1
Xrepeater543 U$$3129/B VGND VGND VPWR VPWR U$$3109/B sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_49_clk _536_/CLK VGND VGND VPWR VPWR _543_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater554 _655_/Q VGND VGND VPWR VPWR U$$2710/B sky130_fd_sc_hd__buf_12
Xrepeater565 U$$2186/B VGND VGND VPWR VPWR U$$2118/B sky130_fd_sc_hd__buf_12
XFILLER_26_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater576 _641_/Q VGND VGND VPWR VPWR U$$1739/B sky130_fd_sc_hd__buf_12
Xrepeater587 U$$1189/B VGND VGND VPWR VPWR U$$1167/B sky130_fd_sc_hd__buf_12
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4280 U$$4280/A U$$4384/A VGND VGND VPWR VPWR U$$4280/X sky130_fd_sc_hd__xor2_1
Xrepeater598 U$$822/A VGND VGND VPWR VPWR U$$778/B sky130_fd_sc_hd__buf_12
XU$$4291 U$$4291/A1 U$$4251/X U$$4291/B1 U$$4252/X VGND VGND VPWR VPWR U$$4292/A sky130_fd_sc_hd__a22o_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3590 U$$28/A1 U$$3624/A2 U$$30/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3591/A sky130_fd_sc_hd__a22o_1
XFILLER_53_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_90_1 dadda_fa_4_90_1/A dadda_fa_4_90_1/B dadda_fa_4_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/B dadda_fa_5_90_1/B sky130_fd_sc_hd__fa_1
XFILLER_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_83_0 dadda_fa_4_83_0/A dadda_fa_4_83_0/B dadda_fa_4_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/A dadda_fa_5_83_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_104_3 dadda_fa_3_104_3/A dadda_fa_3_104_3/B dadda_fa_3_104_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_105_1/B dadda_fa_4_104_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$701 U$$16/A1 U$$689/X U$$975/B1 U$$817/B2 VGND VGND VPWR VPWR U$$702/A sky130_fd_sc_hd__a22o_1
X_662_ _669_/CLK _662_/D VGND VGND VPWR VPWR _662_/Q sky130_fd_sc_hd__dfxtp_1
XU$$712 U$$712/A U$$784/B VGND VGND VPWR VPWR U$$712/X sky130_fd_sc_hd__xor2_1
XU$$723 U$$38/A1 U$$689/X U$$40/A1 U$$817/B2 VGND VGND VPWR VPWR U$$724/A sky130_fd_sc_hd__a22o_1
XFILLER_90_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$734 U$$734/A U$$784/B VGND VGND VPWR VPWR U$$734/X sky130_fd_sc_hd__xor2_1
XU$$745 U$$60/A1 U$$785/A2 U$$62/A1 U$$785/B2 VGND VGND VPWR VPWR U$$746/A sky130_fd_sc_hd__a22o_1
XU$$756 U$$756/A U$$784/B VGND VGND VPWR VPWR U$$756/X sky130_fd_sc_hd__xor2_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_593_ _667_/CLK _593_/D VGND VGND VPWR VPWR _593_/Q sky130_fd_sc_hd__dfxtp_4
XU$$767 U$$82/A1 U$$785/A2 U$$84/A1 U$$785/B2 VGND VGND VPWR VPWR U$$768/A sky130_fd_sc_hd__a22o_1
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$778 U$$778/A U$$778/B VGND VGND VPWR VPWR U$$778/X sky130_fd_sc_hd__xor2_1
XU$$789 U$$926/A1 U$$817/A2 U$$928/A1 U$$817/B2 VGND VGND VPWR VPWR U$$790/A sky130_fd_sc_hd__a22o_1
XFILLER_32_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR _431_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_188_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_98_0 dadda_fa_6_98_0/A dadda_fa_6_98_0/B dadda_fa_6_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_99_0/B dadda_fa_7_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_733__785 VGND VGND VPWR VPWR _733__785/HI U$$2463/B1 sky130_fd_sc_hd__conb_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_40_4 dadda_fa_2_40_4/A dadda_fa_2_40_4/B dadda_fa_2_40_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_1/CIN dadda_fa_3_40_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_33_3 U$$1270/X U$$1403/X U$$1536/X VGND VGND VPWR VPWR dadda_fa_3_34_1/B
+ dadda_fa_3_33_3/B sky130_fd_sc_hd__fa_1
XU$$2130 U$$2130/A U$$2186/B VGND VGND VPWR VPWR U$$2130/X sky130_fd_sc_hd__xor2_1
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2141 U$$908/A1 U$$2161/A2 U$$88/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2142/A sky130_fd_sc_hd__a22o_1
XU$$2152 U$$2152/A _647_/Q VGND VGND VPWR VPWR U$$2152/X sky130_fd_sc_hd__xor2_1
XU$$2163 U$$928/B1 U$$2189/A2 U$$4494/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2164/A
+ sky130_fd_sc_hd__a22o_1
XU$$2174 U$$2174/A U$$2192/A VGND VGND VPWR VPWR U$$2174/X sky130_fd_sc_hd__xor2_1
XU$$1440 U$$892/A1 U$$1472/A2 U$$892/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1441/A sky130_fd_sc_hd__a22o_1
XFILLER_22_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2185 U$$4514/A1 U$$2189/A2 U$$952/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2186/A
+ sky130_fd_sc_hd__a22o_1
XU$$1451 U$$1451/A U$$1505/B VGND VGND VPWR VPWR U$$1451/X sky130_fd_sc_hd__xor2_1
XFILLER_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2196 U$$2194/Y _648_/Q U$$2192/A U$$2195/X U$$2192/Y VGND VGND VPWR VPWR U$$2196/X
+ sky130_fd_sc_hd__a32o_4
XU$$1462 U$$92/A1 U$$1472/A2 U$$94/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1463/A sky130_fd_sc_hd__a22o_1
XU$$1473 U$$1473/A U$$1505/B VGND VGND VPWR VPWR U$$1473/X sky130_fd_sc_hd__xor2_1
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1484 U$$799/A1 U$$1374/X _606_/Q U$$1375/X VGND VGND VPWR VPWR U$$1485/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1495 U$$1495/A _637_/Q VGND VGND VPWR VPWR U$$1495/X sky130_fd_sc_hd__xor2_1
XFILLER_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_78_5 U$$3222/X U$$3355/X U$$3488/X VGND VGND VPWR VPWR dadda_fa_2_79_2/A
+ dadda_fa_2_78_5/A sky130_fd_sc_hd__fa_1
XFILLER_83_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$103 _527_/Q _399_/Q VGND VGND VPWR VPWR final_adder.U$$231/B1 final_adder.U$$725/A
+ sky130_fd_sc_hd__ha_1
XFILLER_170_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$114 _538_/Q _410_/Q VGND VGND VPWR VPWR final_adder.U$$609/B1 final_adder.U$$736/A
+ sky130_fd_sc_hd__ha_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_682__902 VGND VGND VPWR VPWR _682__902/HI _682__902/LO sky130_fd_sc_hd__conb_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$125 _549_/Q _421_/Q VGND VGND VPWR VPWR final_adder.U$$253/B1 final_adder.U$$747/A
+ sky130_fd_sc_hd__ha_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$136 final_adder.U$$9/SUM final_adder.U$$8/SUM VGND VGND VPWR VPWR
+ final_adder.U$$260/B sky130_fd_sc_hd__and2_1
XFILLER_46_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$147 final_adder.U$$641/A final_adder.U$$513/B1 final_adder.U$$147/B1
+ VGND VGND VPWR VPWR final_adder.U$$147/X sky130_fd_sc_hd__a21o_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$158 final_adder.U$$653/A final_adder.U$$652/A VGND VGND VPWR VPWR
+ final_adder.U$$270/A sky130_fd_sc_hd__and2_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$169 final_adder.U$$663/A final_adder.U$$535/B1 final_adder.U$$169/B1
+ VGND VGND VPWR VPWR final_adder.U$$169/X sky130_fd_sc_hd__a21o_1
XFILLER_26_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater395 U$$545/A2 VGND VGND VPWR VPWR U$$491/A2 sky130_fd_sc_hd__buf_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_717__769 VGND VGND VPWR VPWR _717__769/HI U$$1376/A1 sky130_fd_sc_hd__conb_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_102_0 U$$4068/X U$$4201/X U$$4334/X VGND VGND VPWR VPWR dadda_fa_4_103_0/B
+ dadda_fa_4_102_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 b[50] VGND VGND VPWR VPWR _602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 b[60] VGND VGND VPWR VPWR _612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput132 c[102] VGND VGND VPWR VPWR input132/X sky130_fd_sc_hd__clkbuf_4
Xinput143 c[112] VGND VGND VPWR VPWR input143/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_3_50_3 dadda_fa_3_50_3/A dadda_fa_3_50_3/B dadda_fa_3_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/B dadda_fa_4_50_2/CIN sky130_fd_sc_hd__fa_1
Xinput154 c[122] VGND VGND VPWR VPWR input154/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_0_66_3 U$$1336/X U$$1469/X U$$1602/X VGND VGND VPWR VPWR dadda_fa_1_67_6/B
+ dadda_fa_1_66_8/B sky130_fd_sc_hd__fa_1
XFILLER_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput165 c[17] VGND VGND VPWR VPWR input165/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput176 c[27] VGND VGND VPWR VPWR input176/X sky130_fd_sc_hd__buf_2
Xdadda_fa_3_43_2 dadda_fa_3_43_2/A dadda_fa_3_43_2/B dadda_fa_3_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/A dadda_fa_4_43_2/B sky130_fd_sc_hd__fa_1
Xinput187 c[37] VGND VGND VPWR VPWR input187/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput198 c[47] VGND VGND VPWR VPWR input198/X sky130_fd_sc_hd__buf_2
Xdadda_fa_0_59_2 U$$923/X U$$1056/X U$$1189/X VGND VGND VPWR VPWR dadda_fa_1_60_7/A
+ dadda_fa_1_59_8/CIN sky130_fd_sc_hd__fa_2
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$670 final_adder.U$$670/A final_adder.U$$670/B VGND VGND VPWR VPWR
+ _216_/D sky130_fd_sc_hd__xor2_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$681 final_adder.U$$681/A final_adder.U$$681/B VGND VGND VPWR VPWR
+ _227_/D sky130_fd_sc_hd__xor2_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_1 dadda_fa_3_36_1/A dadda_fa_3_36_1/B dadda_fa_3_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/CIN dadda_fa_4_36_2/A sky130_fd_sc_hd__fa_2
XU$$520 U$$520/A U$$547/A VGND VGND VPWR VPWR U$$520/X sky130_fd_sc_hd__xor2_1
X_645_ _645_/CLK _645_/D VGND VGND VPWR VPWR _645_/Q sky130_fd_sc_hd__dfxtp_2
Xfinal_adder.U$$692 final_adder.U$$692/A final_adder.U$$692/B VGND VGND VPWR VPWR
+ _238_/D sky130_fd_sc_hd__xor2_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$531 U$$942/A1 U$$415/X U$$944/A1 U$$416/X VGND VGND VPWR VPWR U$$532/A sky130_fd_sc_hd__a22o_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$542 U$$542/A _623_/Q VGND VGND VPWR VPWR U$$542/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_13_0 dadda_fa_6_13_0/A dadda_fa_6_13_0/B dadda_fa_6_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_14_0/B dadda_fa_7_13_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$553 U$$551/B _623_/Q _624_/Q U$$548/Y VGND VGND VPWR VPWR U$$553/X sky130_fd_sc_hd__a22o_4
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_0 U$$1528/X U$$1661/X U$$1794/X VGND VGND VPWR VPWR dadda_fa_4_30_0/B
+ dadda_fa_4_29_1/CIN sky130_fd_sc_hd__fa_2
XU$$564 U$$16/A1 U$$626/A2 U$$18/A1 U$$553/X VGND VGND VPWR VPWR U$$565/A sky130_fd_sc_hd__a22o_1
XU$$575 U$$575/A U$$623/B VGND VGND VPWR VPWR U$$575/X sky130_fd_sc_hd__xor2_1
XFILLER_45_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_576_ _576_/CLK _576_/D VGND VGND VPWR VPWR _576_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$586 U$$38/A1 U$$626/A2 U$$40/A1 U$$553/X VGND VGND VPWR VPWR U$$587/A sky130_fd_sc_hd__a22o_1
XFILLER_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$597 U$$597/A U$$623/B VGND VGND VPWR VPWR U$$597/X sky130_fd_sc_hd__xor2_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_95_5 input251/X dadda_fa_2_95_5/B dadda_fa_2_95_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_96_2/A dadda_fa_4_95_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_88_4 dadda_fa_2_88_4/A dadda_fa_2_88_4/B dadda_fa_2_88_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/CIN dadda_fa_3_88_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_181_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_25_1 U$$456/X U$$589/X VGND VGND VPWR VPWR dadda_fa_3_26_3/A dadda_fa_4_25_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_707__927 VGND VGND VPWR VPWR _707__927/HI _707__927/LO sky130_fd_sc_hd__conb_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_31_0 U$$69/X U$$202/X U$$335/X VGND VGND VPWR VPWR dadda_fa_3_32_0/CIN
+ dadda_fa_3_31_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1270 U$$1270/A U$$1342/B VGND VGND VPWR VPWR U$$1270/X sky130_fd_sc_hd__xor2_1
XU$$1281 U$$48/A1 U$$1341/A2 U$$50/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1282/A sky130_fd_sc_hd__a22o_1
XU$$1292 U$$1292/A U$$1369/A VGND VGND VPWR VPWR U$$1292/X sky130_fd_sc_hd__xor2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_118_0 dadda_fa_5_118_0/A dadda_fa_5_118_0/B dadda_fa_5_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/A dadda_fa_6_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_83_3 U$$2567/X U$$2700/X U$$2833/X VGND VGND VPWR VPWR dadda_fa_2_84_2/CIN
+ dadda_fa_2_83_5/A sky130_fd_sc_hd__fa_2
XFILLER_85_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_60_2 dadda_fa_4_60_2/A dadda_fa_4_60_2/B dadda_fa_4_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/CIN dadda_fa_5_60_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_76_2 U$$2287/X U$$2420/X U$$2553/X VGND VGND VPWR VPWR dadda_fa_2_77_1/A
+ dadda_fa_2_76_4/A sky130_fd_sc_hd__fa_1
XFILLER_113_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_53_1 dadda_fa_4_53_1/A dadda_fa_4_53_1/B dadda_fa_4_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/B dadda_fa_5_53_1/B sky130_fd_sc_hd__fa_2
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_69_1 U$$2805/X U$$2938/X U$$3071/X VGND VGND VPWR VPWR dadda_fa_2_70_0/CIN
+ dadda_fa_2_69_3/CIN sky130_fd_sc_hd__fa_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_30_0 dadda_fa_7_30_0/A dadda_fa_7_30_0/B dadda_fa_7_30_0/CIN VGND VGND
+ VPWR VPWR _455_/D _326_/D sky130_fd_sc_hd__fa_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_46_0 dadda_fa_4_46_0/A dadda_fa_4_46_0/B dadda_fa_4_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/A dadda_fa_5_46_1/A sky130_fd_sc_hd__fa_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_430_ _432_/CLK _430_/D VGND VGND VPWR VPWR _430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_361_ _367_/CLK _361_/D VGND VGND VPWR VPWR _361_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_292_ _612_/CLK _292_/D VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_98_3 dadda_fa_3_98_3/A dadda_fa_3_98_3/B dadda_fa_3_98_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/B dadda_fa_4_98_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_72_3 U$$1747/X U$$1880/X VGND VGND VPWR VPWR dadda_fa_1_73_8/A dadda_fa_2_72_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_71_1 U$$947/X U$$1080/X U$$1213/X VGND VGND VPWR VPWR dadda_fa_1_72_7/A
+ dadda_fa_1_71_8/B sky130_fd_sc_hd__fa_2
XFILLER_114_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_64_0 U$$135/X U$$268/X U$$401/X VGND VGND VPWR VPWR dadda_fa_1_65_5/B
+ dadda_fa_1_64_7/B sky130_fd_sc_hd__fa_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_845__897 VGND VGND VPWR VPWR _845__897/HI U$$956/B1 sky130_fd_sc_hd__conb_1
XFILLER_91_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$350 U$$759/B1 U$$278/X U$$78/A1 U$$279/X VGND VGND VPWR VPWR U$$351/A sky130_fd_sc_hd__a22o_1
XFILLER_45_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_628_ _633_/CLK _628_/D VGND VGND VPWR VPWR _628_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$361 U$$361/A U$$391/B VGND VGND VPWR VPWR U$$361/X sky130_fd_sc_hd__xor2_1
XFILLER_32_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$372 U$$98/A1 U$$278/X U$$98/B1 U$$279/X VGND VGND VPWR VPWR U$$373/A sky130_fd_sc_hd__a22o_1
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$383 U$$383/A _621_/Q VGND VGND VPWR VPWR U$$383/X sky130_fd_sc_hd__xor2_1
XFILLER_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$394 U$$942/A1 U$$278/X U$$944/A1 U$$279/X VGND VGND VPWR VPWR U$$395/A sky130_fd_sc_hd__a22o_1
X_559_ _633_/CLK _559_/D VGND VGND VPWR VPWR _559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_739__791 VGND VGND VPWR VPWR _739__791/HI U$$2746/A1 sky130_fd_sc_hd__conb_1
XFILLER_173_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_93_2 U$$3651/X U$$3784/X U$$3917/X VGND VGND VPWR VPWR dadda_fa_3_94_1/A
+ dadda_fa_3_93_3/A sky130_fd_sc_hd__fa_1
XFILLER_160_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_70_1 dadda_fa_5_70_1/A dadda_fa_5_70_1/B dadda_fa_5_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/B dadda_fa_7_70_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_86_1 U$$4169/X U$$4302/X U$$4435/X VGND VGND VPWR VPWR dadda_fa_3_87_0/CIN
+ dadda_fa_3_86_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_63_0 dadda_fa_5_63_0/A dadda_fa_5_63_0/B dadda_fa_5_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/A dadda_fa_6_63_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_79_0 dadda_fa_2_79_0/A dadda_fa_2_79_0/B dadda_fa_2_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/B dadda_fa_3_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_62_8 dadda_fa_1_62_8/A dadda_fa_1_62_8/B dadda_fa_1_62_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_3/A dadda_fa_3_62_0/A sky130_fd_sc_hd__fa_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_55_7 U$$3575/X U$$3708/X input207/X VGND VGND VPWR VPWR dadda_fa_2_56_2/CIN
+ dadda_fa_2_55_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_48_6 U$$2497/X U$$2630/X U$$2763/X VGND VGND VPWR VPWR dadda_fa_2_49_3/A
+ dadda_fa_2_48_5/CIN sky130_fd_sc_hd__fa_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_78_0 dadda_fa_7_78_0/A dadda_fa_7_78_0/B dadda_fa_7_78_0/CIN VGND VGND
+ VPWR VPWR _503_/D _374_/D sky130_fd_sc_hd__fa_1
XFILLER_163_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_81_0 U$$1232/Y U$$1366/X U$$1499/X VGND VGND VPWR VPWR dadda_fa_2_82_1/A
+ dadda_fa_2_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4109 U$$4109/A VGND VGND VPWR VPWR U$$4109/Y sky130_fd_sc_hd__inv_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3408 U$$4504/A1 U$$3292/X U$$4506/A1 U$$3293/X VGND VGND VPWR VPWR U$$3409/A sky130_fd_sc_hd__a22o_1
XFILLER_86_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3419 U$$3419/A _665_/Q VGND VGND VPWR VPWR U$$3419/X sky130_fd_sc_hd__xor2_1
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2707 U$$787/B1 U$$2729/A2 U$$654/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2708/A sky130_fd_sc_hd__a22o_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2718 U$$2718/A _655_/Q VGND VGND VPWR VPWR U$$2718/X sky130_fd_sc_hd__xor2_1
XFILLER_27_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2729 U$$4510/A1 U$$2729/A2 U$$950/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2730/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _601_/CLK _413_/D VGND VGND VPWR VPWR _413_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _480_/CLK _344_/D VGND VGND VPWR VPWR _344_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_275_ _280_/CLK _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_80_0 dadda_fa_6_80_0/A dadda_fa_6_80_0/B dadda_fa_6_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_81_0/B dadda_fa_7_80_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_96_0 dadda_fa_3_96_0/A dadda_fa_3_96_0/B dadda_fa_3_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/B dadda_fa_4_96_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_143_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_58_5 dadda_fa_2_58_5/A dadda_fa_2_58_5/B dadda_fa_2_58_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_2/A dadda_fa_4_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3920 _590_/Q U$$3840/X _591_/Q U$$3841/X VGND VGND VPWR VPWR U$$3921/A sky130_fd_sc_hd__a22o_1
XFILLER_76_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3931 U$$3931/A _673_/Q VGND VGND VPWR VPWR U$$3931/X sky130_fd_sc_hd__xor2_1
XU$$3942 U$$654/A1 U$$3970/A2 U$$4492/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3943/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3953 U$$3953/A _673_/Q VGND VGND VPWR VPWR U$$3953/X sky130_fd_sc_hd__xor2_1
XFILLER_92_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3964 U$$539/A1 U$$3970/A2 _613_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3965/A sky130_fd_sc_hd__a22o_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3975 U$$4058/B VGND VGND VPWR VPWR U$$3975/Y sky130_fd_sc_hd__inv_1
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3986 U$$3986/A U$$4044/B VGND VGND VPWR VPWR U$$3986/X sky130_fd_sc_hd__xor2_1
XFILLER_64_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3997 U$$4271/A1 U$$4045/A2 U$$4273/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$3998/A
+ sky130_fd_sc_hd__a22o_1
XU$$180 U$$180/A U$$262/B VGND VGND VPWR VPWR U$$180/X sky130_fd_sc_hd__xor2_1
XU$$191 U$$54/A1 U$$141/X U$$56/A1 U$$142/X VGND VGND VPWR VPWR U$$192/A sky130_fd_sc_hd__a22o_1
XFILLER_178_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput266 _276_/Q VGND VGND VPWR VPWR o[108] sky130_fd_sc_hd__buf_2
Xoutput277 _286_/Q VGND VGND VPWR VPWR o[118] sky130_fd_sc_hd__buf_2
Xoutput288 _180_/Q VGND VGND VPWR VPWR o[12] sky130_fd_sc_hd__buf_2
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput299 _190_/Q VGND VGND VPWR VPWR o[22] sky130_fd_sc_hd__buf_2
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_5 U$$3984/X U$$4117/X _677_/Q VGND VGND VPWR VPWR dadda_fa_2_61_2/A
+ dadda_fa_2_60_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_53_4 U$$1975/X U$$2108/X U$$2241/X VGND VGND VPWR VPWR dadda_fa_2_54_1/CIN
+ dadda_fa_2_53_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_46_3 U$$1296/X U$$1429/X U$$1562/X VGND VGND VPWR VPWR dadda_fa_2_47_2/CIN
+ dadda_fa_2_46_5/A sky130_fd_sc_hd__fa_2
XFILLER_55_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_23_2 dadda_fa_4_23_2/A dadda_fa_4_23_2/B dadda_fa_4_23_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/CIN dadda_fa_5_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_16_1 U$$1103/X U$$1189/B input164/X VGND VGND VPWR VPWR dadda_fa_5_17_0/B
+ dadda_fa_5_16_1/B sky130_fd_sc_hd__fa_1
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3205 U$$4438/A1 U$$3243/A2 U$$4303/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3206/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3216 U$$3216/A U$$3224/B VGND VGND VPWR VPWR U$$3216/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3227 U$$76/A1 U$$3243/A2 U$$76/B1 U$$3243/B2 VGND VGND VPWR VPWR U$$3228/A sky130_fd_sc_hd__a22o_1
XFILLER_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3238 U$$3238/A _663_/Q VGND VGND VPWR VPWR U$$3238/X sky130_fd_sc_hd__xor2_1
XU$$2504 U$$4285/A1 U$$2534/A2 U$$3191/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2505/A
+ sky130_fd_sc_hd__a22o_1
XU$$3249 _597_/Q U$$3155/X _598_/Q U$$3156/X VGND VGND VPWR VPWR U$$3250/A sky130_fd_sc_hd__a22o_1
XFILLER_19_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2515 U$$2515/A U$$2585/B VGND VGND VPWR VPWR U$$2515/X sky130_fd_sc_hd__xor2_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2526 _578_/Q U$$2534/A2 U$$4446/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2527/A sky130_fd_sc_hd__a22o_1
XFILLER_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2537 U$$2537/A U$$2585/B VGND VGND VPWR VPWR U$$2537/X sky130_fd_sc_hd__xor2_1
XU$$2548 _589_/Q U$$2470/X _590_/Q U$$2471/X VGND VGND VPWR VPWR U$$2549/A sky130_fd_sc_hd__a22o_1
XU$$1803 U$$979/B1 U$$1903/A2 U$$4271/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1804/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2559 U$$2559/A _653_/Q VGND VGND VPWR VPWR U$$2559/X sky130_fd_sc_hd__xor2_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1814 U$$1814/A U$$1918/A VGND VGND VPWR VPWR U$$1814/X sky130_fd_sc_hd__xor2_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1825 U$$4291/A1 U$$1897/A2 U$$868/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1826/A
+ sky130_fd_sc_hd__a22o_1
XU$$1836 U$$1836/A U$$1918/A VGND VGND VPWR VPWR U$$1836/X sky130_fd_sc_hd__xor2_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1847 U$$3489/B1 U$$1903/A2 U$$3217/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1848/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1858 U$$1858/A U$$1918/A VGND VGND VPWR VPWR U$$1858/X sky130_fd_sc_hd__xor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1869 U$$88/A1 U$$1897/A2 U$$912/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1870/A sky130_fd_sc_hd__a22o_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_327_ _327_/CLK _327_/D VGND VGND VPWR VPWR _327_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_258_ _503_/CLK _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_189_ _329_/CLK _189_/D VGND VGND VPWR VPWR _189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_70_4 dadda_fa_2_70_4/A dadda_fa_2_70_4/B dadda_fa_2_70_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/CIN dadda_fa_3_70_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_63_3 dadda_fa_2_63_3/A dadda_fa_2_63_3/B dadda_fa_2_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/B dadda_fa_3_63_3/B sky130_fd_sc_hd__fa_1
XFILLER_111_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater703 _577_/Q VGND VGND VPWR VPWR U$$4442/A1 sky130_fd_sc_hd__buf_12
XFILLER_111_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater714 _573_/Q VGND VGND VPWR VPWR U$$735/A1 sky130_fd_sc_hd__buf_12
XFILLER_78_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater725 U$$4424/A1 VGND VGND VPWR VPWR U$$40/A1 sky130_fd_sc_hd__buf_12
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_56_2 dadda_fa_2_56_2/A dadda_fa_2_56_2/B dadda_fa_2_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/A dadda_fa_3_56_3/A sky130_fd_sc_hd__fa_2
Xrepeater736 _563_/Q VGND VGND VPWR VPWR U$$30/A1 sky130_fd_sc_hd__buf_12
Xrepeater747 _558_/Q VGND VGND VPWR VPWR U$$842/A1 sky130_fd_sc_hd__buf_12
Xrepeater758 U$$969/A1 VGND VGND VPWR VPWR U$$8/B1 sky130_fd_sc_hd__buf_12
XFILLER_77_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4440 _576_/Q U$$4388/X U$$4442/A1 U$$4389/X VGND VGND VPWR VPWR U$$4441/A sky130_fd_sc_hd__a22o_2
XFILLER_37_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_33_1 dadda_fa_5_33_1/A dadda_fa_5_33_1/B dadda_fa_5_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/B dadda_fa_7_33_0/A sky130_fd_sc_hd__fa_1
XU$$4451 U$$4451/A U$$4451/B VGND VGND VPWR VPWR U$$4451/X sky130_fd_sc_hd__xor2_1
XU$$4462 U$$78/A1 U$$4388/X U$$765/A1 U$$4389/X VGND VGND VPWR VPWR U$$4463/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_1 dadda_fa_2_49_1/A dadda_fa_2_49_1/B dadda_fa_2_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_0/CIN dadda_fa_3_49_2/CIN sky130_fd_sc_hd__fa_1
XU$$4473 U$$4473/A U$$4473/B VGND VGND VPWR VPWR U$$4473/X sky130_fd_sc_hd__xor2_1
XU$$4484 U$$4484/A1 U$$4388/X U$$4486/A1 U$$4389/X VGND VGND VPWR VPWR U$$4485/A sky130_fd_sc_hd__a22o_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3750 U$$3750/A U$$3784/B VGND VGND VPWR VPWR U$$3750/X sky130_fd_sc_hd__xor2_1
XFILLER_53_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_26_0 dadda_fa_5_26_0/A dadda_fa_5_26_0/B dadda_fa_5_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/A dadda_fa_6_26_0/CIN sky130_fd_sc_hd__fa_1
XU$$4495 U$$4495/A U$$4495/B VGND VGND VPWR VPWR U$$4495/X sky130_fd_sc_hd__xor2_1
XFILLER_53_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3761 U$$4446/A1 U$$3795/A2 _580_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3762/A sky130_fd_sc_hd__a22o_1
XU$$3772 U$$3772/A U$$3794/B VGND VGND VPWR VPWR U$$3772/X sky130_fd_sc_hd__xor2_1
XU$$3783 U$$632/A1 U$$3783/A2 U$$771/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3784/A sky130_fd_sc_hd__a22o_1
XFILLER_53_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3794 U$$3794/A U$$3794/B VGND VGND VPWR VPWR U$$3794/X sky130_fd_sc_hd__xor2_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_100_0 dadda_fa_5_100_0/A dadda_fa_5_100_0/B dadda_fa_5_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/A dadda_fa_6_100_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_51_1 U$$508/X U$$641/X U$$774/X VGND VGND VPWR VPWR dadda_fa_2_52_0/CIN
+ dadda_fa_2_51_3/CIN sky130_fd_sc_hd__fa_1
XU$$905 U$$905/A U$$923/B VGND VGND VPWR VPWR U$$905/X sky130_fd_sc_hd__xor2_1
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$916 U$$92/B1 U$$928/A2 U$$96/A1 U$$928/B2 VGND VGND VPWR VPWR U$$917/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_0 U$$95/X U$$228/X U$$361/X VGND VGND VPWR VPWR dadda_fa_2_45_2/B dadda_fa_2_44_4/B
+ sky130_fd_sc_hd__fa_2
XU$$927 U$$927/A U$$943/B VGND VGND VPWR VPWR U$$927/X sky130_fd_sc_hd__xor2_1
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$938 U$$938/A1 U$$826/X _607_/Q U$$827/X VGND VGND VPWR VPWR U$$939/A sky130_fd_sc_hd__a22o_1
XU$$949 U$$949/A _629_/Q VGND VGND VPWR VPWR U$$949/X sky130_fd_sc_hd__xor2_1
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_3 dadda_fa_3_80_3/A dadda_fa_3_80_3/B dadda_fa_3_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/B dadda_fa_4_80_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_166_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_73_2 dadda_fa_3_73_2/A dadda_fa_3_73_2/B dadda_fa_3_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/A dadda_fa_4_73_2/B sky130_fd_sc_hd__fa_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_66_1 dadda_fa_3_66_1/A dadda_fa_3_66_1/B dadda_fa_3_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/CIN dadda_fa_4_66_2/A sky130_fd_sc_hd__fa_1
XFILLER_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_43_0 dadda_fa_6_43_0/A dadda_fa_6_43_0/B dadda_fa_6_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_44_0/B dadda_fa_7_43_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_59_0 dadda_fa_3_59_0/A dadda_fa_3_59_0/B dadda_fa_3_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/B dadda_fa_4_59_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3002 U$$3002/A U$$3004/B VGND VGND VPWR VPWR U$$3002/X sky130_fd_sc_hd__xor2_1
XU$$3013 _659_/Q VGND VGND VPWR VPWR U$$3013/Y sky130_fd_sc_hd__inv_1
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3024 _553_/Q U$$3090/A2 U$$4122/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3025/A sky130_fd_sc_hd__a22o_1
XU$$3035 U$$3035/A U$$3085/B VGND VGND VPWR VPWR U$$3035/X sky130_fd_sc_hd__xor2_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3046 _564_/Q U$$3090/A2 _565_/Q U$$3090/B2 VGND VGND VPWR VPWR U$$3047/A sky130_fd_sc_hd__a22o_1
XU$$2301 U$$2301/A U$$2327/B VGND VGND VPWR VPWR U$$2301/X sky130_fd_sc_hd__xor2_1
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2312 U$$942/A1 U$$2326/A2 U$$4506/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2313/A
+ sky130_fd_sc_hd__a22o_1
XU$$3057 U$$3057/A U$$3085/B VGND VGND VPWR VPWR U$$3057/X sky130_fd_sc_hd__xor2_1
XFILLER_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2323 U$$2323/A _649_/Q VGND VGND VPWR VPWR U$$2323/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_2 dadda_fa_4_102_2/A dadda_fa_4_102_2/B dadda_fa_4_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/CIN dadda_fa_5_102_1/CIN sky130_fd_sc_hd__fa_1
XU$$3068 U$$876/A1 U$$3090/A2 U$$4303/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3069/A
+ sky130_fd_sc_hd__a22o_1
XU$$2334 U$$2332/B _649_/Q _650_/Q U$$2329/Y VGND VGND VPWR VPWR U$$2334/X sky130_fd_sc_hd__a22o_4
XU$$3079 U$$3079/A U$$3137/B VGND VGND VPWR VPWR U$$3079/X sky130_fd_sc_hd__xor2_1
XU$$1600 U$$1600/A _639_/Q VGND VGND VPWR VPWR U$$1600/X sky130_fd_sc_hd__xor2_1
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2345 U$$16/A1 U$$2333/X U$$18/A1 U$$2334/X VGND VGND VPWR VPWR U$$2346/A sky130_fd_sc_hd__a22o_1
XU$$2356 U$$2356/A U$$2436/B VGND VGND VPWR VPWR U$$2356/X sky130_fd_sc_hd__xor2_1
XU$$1611 U$$787/B1 U$$1641/A2 U$$654/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1612/A sky130_fd_sc_hd__a22o_1
XU$$2367 U$$4285/A1 U$$2421/A2 U$$3191/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2368/A
+ sky130_fd_sc_hd__a22o_1
XU$$1622 U$$1622/A _639_/Q VGND VGND VPWR VPWR U$$1622/X sky130_fd_sc_hd__xor2_1
XU$$2378 U$$2378/A U$$2436/B VGND VGND VPWR VPWR U$$2378/X sky130_fd_sc_hd__xor2_1
XU$$1633 U$$948/A1 U$$1641/A2 U$$950/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1634/A sky130_fd_sc_hd__a22o_1
XU$$1644 _639_/Q VGND VGND VPWR VPWR U$$1644/Y sky130_fd_sc_hd__inv_1
XU$$2389 _578_/Q U$$2421/A2 U$$4446/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2390/A sky130_fd_sc_hd__a22o_1
XU$$1655 U$$1655/A U$$1727/B VGND VGND VPWR VPWR U$$1655/X sky130_fd_sc_hd__xor2_1
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1666 U$$979/B1 U$$1734/A2 U$$983/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1667/A sky130_fd_sc_hd__a22o_1
XFILLER_188_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1677 U$$1677/A U$$1781/A VGND VGND VPWR VPWR U$$1677/X sky130_fd_sc_hd__xor2_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1688 U$$4291/A1 U$$1726/A2 U$$868/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1689/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1699 U$$1699/A U$$1727/B VGND VGND VPWR VPWR U$$1699/X sky130_fd_sc_hd__xor2_1
XFILLER_30_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_116_0 dadda_fa_7_116_0/A dadda_fa_7_116_0/B dadda_fa_7_116_0/CIN VGND
+ VGND VPWR VPWR _541_/D _412_/D sky130_fd_sc_hd__fa_2
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_0 dadda_fa_2_61_0/A dadda_fa_2_61_0/B dadda_fa_2_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/B dadda_fa_3_61_2/B sky130_fd_sc_hd__fa_1
Xrepeater500 U$$1897/B2 VGND VGND VPWR VPWR U$$1903/B2 sky130_fd_sc_hd__buf_12
XFILLER_112_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$307 final_adder.U$$306/A final_adder.U$$229/X final_adder.U$$231/X
+ VGND VGND VPWR VPWR final_adder.U$$307/X sky130_fd_sc_hd__a21o_1
Xrepeater511 U$$1238/X VGND VGND VPWR VPWR U$$1341/B2 sky130_fd_sc_hd__buf_12
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater522 _675_/Q VGND VGND VPWR VPWR U$$4058/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$329 final_adder.U$$328/A final_adder.U$$273/X final_adder.U$$275/X
+ VGND VGND VPWR VPWR final_adder.U$$329/X sky130_fd_sc_hd__a21o_1
Xrepeater533 _667_/Q VGND VGND VPWR VPWR U$$3561/A sky130_fd_sc_hd__buf_12
XFILLER_38_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater544 U$$3137/B VGND VGND VPWR VPWR U$$3129/B sky130_fd_sc_hd__buf_12
Xrepeater555 _653_/Q VGND VGND VPWR VPWR U$$2533/B sky130_fd_sc_hd__buf_12
Xrepeater566 _647_/Q VGND VGND VPWR VPWR U$$2186/B sky130_fd_sc_hd__buf_12
Xrepeater577 _641_/Q VGND VGND VPWR VPWR U$$1781/A sky130_fd_sc_hd__buf_12
Xrepeater588 _633_/Q VGND VGND VPWR VPWR U$$1189/B sky130_fd_sc_hd__buf_12
XFILLER_168_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4270 U$$4270/A U$$4384/A VGND VGND VPWR VPWR U$$4270/X sky130_fd_sc_hd__xor2_1
XFILLER_53_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4281 _565_/Q U$$4377/A2 _566_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4282/A sky130_fd_sc_hd__a22o_1
Xrepeater599 _627_/Q VGND VGND VPWR VPWR U$$822/A sky130_fd_sc_hd__buf_12
XU$$4292 U$$4292/A U$$4332/B VGND VGND VPWR VPWR U$$4292/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3580 U$$4265/A1 U$$3624/A2 U$$979/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3581/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3591 U$$3591/A U$$3625/B VGND VGND VPWR VPWR U$$3591/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2890 U$$2890/A U$$2996/B VGND VGND VPWR VPWR U$$2890/X sky130_fd_sc_hd__xor2_1
XFILLER_139_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_90_2 dadda_fa_4_90_2/A dadda_fa_4_90_2/B dadda_fa_4_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/CIN dadda_fa_5_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_83_1 dadda_fa_4_83_1/A dadda_fa_4_83_1/B dadda_fa_4_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/B dadda_fa_5_83_1/B sky130_fd_sc_hd__fa_1
XFILLER_162_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_60_0 dadda_fa_7_60_0/A dadda_fa_7_60_0/B dadda_fa_7_60_0/CIN VGND VGND
+ VPWR VPWR _485_/D _356_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_76_0 dadda_fa_4_76_0/A dadda_fa_4_76_0/B dadda_fa_4_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/A dadda_fa_5_76_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_661_ _669_/CLK _661_/D VGND VGND VPWR VPWR _661_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$702 U$$702/A U$$784/B VGND VGND VPWR VPWR U$$702/X sky130_fd_sc_hd__xor2_1
XFILLER_152_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$713 U$$987/A1 U$$785/A2 U$$28/B1 U$$785/B2 VGND VGND VPWR VPWR U$$714/A sky130_fd_sc_hd__a22o_1
XU$$724 U$$724/A U$$784/B VGND VGND VPWR VPWR U$$724/X sky130_fd_sc_hd__xor2_1
XU$$735 U$$735/A1 U$$689/X U$$52/A1 U$$817/B2 VGND VGND VPWR VPWR U$$736/A sky130_fd_sc_hd__a22o_1
XFILLER_72_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_592_ _679_/CLK _592_/D VGND VGND VPWR VPWR _592_/Q sky130_fd_sc_hd__dfxtp_1
XU$$746 U$$746/A U$$778/B VGND VGND VPWR VPWR U$$746/X sky130_fd_sc_hd__xor2_2
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$757 U$$72/A1 U$$785/A2 U$$74/A1 U$$785/B2 VGND VGND VPWR VPWR U$$758/A sky130_fd_sc_hd__a22o_1
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$768 U$$768/A U$$778/B VGND VGND VPWR VPWR U$$768/X sky130_fd_sc_hd__xor2_1
XFILLER_44_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$779 U$$92/B1 U$$785/A2 U$$96/A1 U$$785/B2 VGND VGND VPWR VPWR U$$780/A sky130_fd_sc_hd__a22o_1
XFILLER_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_40_5 dadda_fa_2_40_5/A dadda_fa_2_40_5/B dadda_fa_2_40_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_2/A dadda_fa_4_40_0/A sky130_fd_sc_hd__fa_2
XFILLER_82_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_33_4 U$$1669/X U$$1802/X U$$1935/X VGND VGND VPWR VPWR dadda_fa_3_34_1/CIN
+ dadda_fa_3_33_3/CIN sky130_fd_sc_hd__fa_1
XU$$2120 U$$2120/A _647_/Q VGND VGND VPWR VPWR U$$2120/X sky130_fd_sc_hd__xor2_1
XFILLER_74_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2131 U$$759/B1 U$$2059/X U$$78/A1 U$$2060/X VGND VGND VPWR VPWR U$$2132/A sky130_fd_sc_hd__a22o_1
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2142 U$$2142/A _647_/Q VGND VGND VPWR VPWR U$$2142/X sky130_fd_sc_hd__xor2_1
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2153 U$$98/A1 U$$2189/A2 U$$98/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2154/A sky130_fd_sc_hd__a22o_1
XFILLER_23_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2164 U$$2164/A U$$2192/A VGND VGND VPWR VPWR U$$2164/X sky130_fd_sc_hd__xor2_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2175 U$$942/A1 U$$2189/A2 U$$944/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2176/A sky130_fd_sc_hd__a22o_1
XU$$1430 U$$60/A1 U$$1472/A2 U$$62/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1431/A sky130_fd_sc_hd__a22o_1
XU$$1441 U$$1441/A U$$1505/B VGND VGND VPWR VPWR U$$1441/X sky130_fd_sc_hd__xor2_1
XFILLER_16_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2186 U$$2186/A U$$2186/B VGND VGND VPWR VPWR U$$2186/X sky130_fd_sc_hd__xor2_1
XU$$2197 U$$2195/B U$$2192/A _648_/Q U$$2192/Y VGND VGND VPWR VPWR U$$2197/X sky130_fd_sc_hd__a22o_4
XU$$1452 U$$902/B1 U$$1472/A2 U$$84/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1453/A sky130_fd_sc_hd__a22o_1
XU$$1463 U$$1463/A U$$1479/B VGND VGND VPWR VPWR U$$1463/X sky130_fd_sc_hd__xor2_1
XU$$1474 U$$787/B1 U$$1474/A2 U$$654/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1475/A sky130_fd_sc_hd__a22o_1
XU$$1485 U$$1485/A U$$1505/B VGND VGND VPWR VPWR U$$1485/X sky130_fd_sc_hd__xor2_1
XU$$1496 U$$948/A1 U$$1374/X U$$950/A1 U$$1375/X VGND VGND VPWR VPWR U$$1497/A sky130_fd_sc_hd__a22o_1
XFILLER_31_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_93_0 dadda_fa_5_93_0/A dadda_fa_5_93_0/B dadda_fa_5_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/A dadda_fa_6_93_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_159_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_78_6 U$$3621/X U$$3754/X U$$3887/X VGND VGND VPWR VPWR dadda_fa_2_79_2/B
+ dadda_fa_2_78_5/B sky130_fd_sc_hd__fa_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$104 _528_/Q _400_/Q VGND VGND VPWR VPWR final_adder.U$$599/B1 final_adder.U$$726/A
+ sky130_fd_sc_hd__ha_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$115 _539_/Q _411_/Q VGND VGND VPWR VPWR final_adder.U$$243/B1 final_adder.U$$737/A
+ sky130_fd_sc_hd__ha_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$126 _550_/Q _422_/Q VGND VGND VPWR VPWR final_adder.U$$621/B1 final_adder.U$$748/A
+ sky130_fd_sc_hd__ha_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$137 final_adder.U$$9/SUM final_adder.U$$8/COUT final_adder.U$$9/COUT
+ VGND VGND VPWR VPWR final_adder.U$$137/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$148 final_adder.U$$643/A final_adder.U$$642/A VGND VGND VPWR VPWR
+ final_adder.U$$266/B sky130_fd_sc_hd__and2_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$159 final_adder.U$$653/A final_adder.U$$525/B1 final_adder.U$$159/B1
+ VGND VGND VPWR VPWR final_adder.U$$159/X sky130_fd_sc_hd__a21o_1
Xrepeater385 U$$1093/A2 VGND VGND VPWR VPWR U$$999/A2 sky130_fd_sc_hd__buf_12
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater396 U$$415/X VGND VGND VPWR VPWR U$$545/A2 sky130_fd_sc_hd__buf_12
XFILLER_54_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_102_1 U$$4467/X input132/X dadda_fa_3_102_1/CIN VGND VGND VPWR VPWR dadda_fa_4_103_0/CIN
+ dadda_fa_4_102_2/A sky130_fd_sc_hd__fa_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 b[41] VGND VGND VPWR VPWR _593_/D sky130_fd_sc_hd__clkbuf_4
Xinput111 b[51] VGND VGND VPWR VPWR _603_/D sky130_fd_sc_hd__clkbuf_1
Xinput122 b[61] VGND VGND VPWR VPWR _613_/D sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_6_123_0 dadda_fa_6_123_0/A dadda_fa_6_123_0/B dadda_fa_6_123_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_124_0/B dadda_fa_7_123_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput133 c[103] VGND VGND VPWR VPWR input133/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput144 c[113] VGND VGND VPWR VPWR input144/X sky130_fd_sc_hd__clkbuf_2
Xinput155 c[123] VGND VGND VPWR VPWR input155/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_0_66_4 U$$1735/X U$$1868/X U$$2001/X VGND VGND VPWR VPWR dadda_fa_1_67_6/CIN
+ dadda_fa_1_66_8/CIN sky130_fd_sc_hd__fa_1
Xinput166 c[18] VGND VGND VPWR VPWR input166/X sky130_fd_sc_hd__clkbuf_2
Xinput177 c[28] VGND VGND VPWR VPWR input177/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_3_43_3 dadda_fa_3_43_3/A dadda_fa_3_43_3/B dadda_fa_3_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/B dadda_fa_4_43_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 c[38] VGND VGND VPWR VPWR input188/X sky130_fd_sc_hd__buf_2
Xinput199 c[48] VGND VGND VPWR VPWR input199/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$660 final_adder.U$$660/A final_adder.U$$660/B VGND VGND VPWR VPWR
+ _206_/D sky130_fd_sc_hd__xor2_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$671 final_adder.U$$671/A final_adder.U$$671/B VGND VGND VPWR VPWR
+ _217_/D sky130_fd_sc_hd__xor2_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_644_ _644_/CLK _644_/D VGND VGND VPWR VPWR _644_/Q sky130_fd_sc_hd__dfxtp_2
XU$$510 U$$510/A U$$547/A VGND VGND VPWR VPWR U$$510/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$682 final_adder.U$$682/A final_adder.U$$682/B VGND VGND VPWR VPWR
+ _228_/D sky130_fd_sc_hd__xor2_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$521 U$$932/A1 U$$545/A2 U$$934/A1 U$$416/X VGND VGND VPWR VPWR U$$522/A sky130_fd_sc_hd__a22o_1
XFILLER_57_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_36_2 dadda_fa_3_36_2/A dadda_fa_3_36_2/B dadda_fa_3_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/A dadda_fa_4_36_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$693 final_adder.U$$693/A final_adder.U$$693/B VGND VGND VPWR VPWR
+ _239_/D sky130_fd_sc_hd__xor2_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$532 U$$532/A _623_/Q VGND VGND VPWR VPWR U$$532/X sky130_fd_sc_hd__xor2_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$543 U$$952/B1 U$$545/A2 U$$956/A1 U$$416/X VGND VGND VPWR VPWR U$$544/A sky130_fd_sc_hd__a22o_1
XFILLER_45_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_29_1 U$$1927/X input178/X dadda_fa_3_29_1/CIN VGND VGND VPWR VPWR dadda_fa_4_30_0/CIN
+ dadda_fa_4_29_2/A sky130_fd_sc_hd__fa_2
XU$$554 U$$554/A1 U$$626/A2 U$$8/A1 U$$553/X VGND VGND VPWR VPWR U$$555/A sky130_fd_sc_hd__a22o_1
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$565 U$$565/A U$$623/B VGND VGND VPWR VPWR U$$565/X sky130_fd_sc_hd__xor2_1
X_575_ _579_/CLK _575_/D VGND VGND VPWR VPWR _575_/Q sky130_fd_sc_hd__dfxtp_4
XU$$576 U$$987/A1 U$$626/A2 U$$28/B1 U$$553/X VGND VGND VPWR VPWR U$$577/A sky130_fd_sc_hd__a22o_1
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$587 U$$587/A U$$623/B VGND VGND VPWR VPWR U$$587/X sky130_fd_sc_hd__xor2_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$598 U$$735/A1 U$$626/A2 U$$52/A1 U$$553/X VGND VGND VPWR VPWR U$$599/A sky130_fd_sc_hd__a22o_1
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_88_5 dadda_fa_2_88_5/A dadda_fa_2_88_5/B dadda_fa_2_88_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_2/A dadda_fa_4_88_0/A sky130_fd_sc_hd__fa_2
XFILLER_141_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_31_1 U$$468/X U$$601/X U$$734/X VGND VGND VPWR VPWR dadda_fa_3_32_1/A
+ dadda_fa_3_31_3/A sky130_fd_sc_hd__fa_2
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_24_0 U$$55/X U$$188/X U$$321/X VGND VGND VPWR VPWR dadda_fa_3_25_3/A dadda_fa_3_24_3/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_168_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1260 U$$1260/A U$$1342/B VGND VGND VPWR VPWR U$$1260/X sky130_fd_sc_hd__xor2_1
XU$$1271 U$$4285/A1 U$$1341/A2 U$$3191/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1282 U$$1282/A U$$1342/B VGND VGND VPWR VPWR U$$1282/X sky130_fd_sc_hd__xor2_1
XU$$1293 U$$60/A1 U$$1341/A2 U$$4446/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1294/A sky130_fd_sc_hd__a22o_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_118_1 dadda_fa_5_118_1/A dadda_fa_5_118_1/B dadda_ha_4_118_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/B dadda_fa_7_118_0/A sky130_fd_sc_hd__fa_1
Xdadda_ha_1_84_6 U$$3766/X U$$3899/X VGND VGND VPWR VPWR dadda_fa_2_85_4/A dadda_fa_3_84_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_176_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_83_4 U$$2966/X U$$3099/X U$$3232/X VGND VGND VPWR VPWR dadda_fa_2_84_3/A
+ dadda_fa_2_83_5/B sky130_fd_sc_hd__fa_2
XFILLER_132_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_76_3 U$$2686/X U$$2819/X U$$2952/X VGND VGND VPWR VPWR dadda_fa_2_77_1/B
+ dadda_fa_2_76_4/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_53_2 dadda_fa_4_53_2/A dadda_fa_4_53_2/B dadda_fa_4_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/CIN dadda_fa_5_53_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_69_2 U$$3204/X U$$3337/X U$$3470/X VGND VGND VPWR VPWR dadda_fa_2_70_1/A
+ dadda_fa_2_69_4/A sky130_fd_sc_hd__fa_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_1 dadda_fa_4_46_1/A dadda_fa_4_46_1/B dadda_fa_4_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/B dadda_fa_5_46_1/B sky130_fd_sc_hd__fa_1
XFILLER_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_23_0 dadda_fa_7_23_0/A dadda_fa_7_23_0/B dadda_fa_7_23_0/CIN VGND VGND
+ VPWR VPWR _448_/D _319_/D sky130_fd_sc_hd__fa_2
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_0 dadda_fa_4_39_0/A dadda_fa_4_39_0/B dadda_fa_4_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/A dadda_fa_5_39_1/A sky130_fd_sc_hd__fa_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _632_/CLK _360_/D VGND VGND VPWR VPWR _360_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_291_ _612_/CLK _291_/D VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_689__909 VGND VGND VPWR VPWR _689__909/HI _689__909/LO sky130_fd_sc_hd__conb_1
XFILLER_1_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_71_2 U$$1346/X U$$1479/X U$$1612/X VGND VGND VPWR VPWR dadda_fa_1_72_7/B
+ dadda_fa_1_71_8/CIN sky130_fd_sc_hd__fa_2
XFILLER_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_64_1 U$$534/X U$$667/X U$$800/X VGND VGND VPWR VPWR dadda_fa_1_65_5/CIN
+ dadda_fa_1_64_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_41_0 dadda_fa_3_41_0/A dadda_fa_3_41_0/B dadda_fa_3_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/B dadda_fa_4_41_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_57_0 U$$121/X U$$254/X U$$387/X VGND VGND VPWR VPWR dadda_fa_1_58_7/A
+ dadda_fa_1_57_8/B sky130_fd_sc_hd__fa_2
XFILLER_114_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_627_ _633_/CLK _627_/D VGND VGND VPWR VPWR _627_/Q sky130_fd_sc_hd__dfxtp_4
XU$$340 U$$66/A1 U$$278/X U$$68/A1 U$$279/X VGND VGND VPWR VPWR U$$341/A sky130_fd_sc_hd__a22o_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$351 U$$351/A U$$357/B VGND VGND VPWR VPWR U$$351/X sky130_fd_sc_hd__xor2_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$362 U$$88/A1 U$$278/X U$$90/A1 U$$279/X VGND VGND VPWR VPWR U$$363/A sky130_fd_sc_hd__a22o_1
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$373 U$$373/A _621_/Q VGND VGND VPWR VPWR U$$373/X sky130_fd_sc_hd__xor2_1
XFILLER_33_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$384 U$$932/A1 U$$278/X U$$934/A1 U$$279/X VGND VGND VPWR VPWR U$$385/A sky130_fd_sc_hd__a22o_1
XFILLER_44_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$395 U$$395/A _621_/Q VGND VGND VPWR VPWR U$$395/X sky130_fd_sc_hd__xor2_1
X_558_ _649_/CLK _558_/D VGND VGND VPWR VPWR _558_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_489_ _490_/CLK _489_/D VGND VGND VPWR VPWR _489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_93_3 U$$4050/X U$$4183/X U$$4316/X VGND VGND VPWR VPWR dadda_fa_3_94_1/B
+ dadda_fa_3_93_3/B sky130_fd_sc_hd__fa_2
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_86_2 input241/X dadda_fa_2_86_2/B dadda_fa_2_86_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_87_1/A dadda_fa_3_86_3/A sky130_fd_sc_hd__fa_2
XFILLER_5_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_63_1 dadda_fa_5_63_1/A dadda_fa_5_63_1/B dadda_fa_5_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/B dadda_fa_7_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_113_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_79_1 dadda_fa_2_79_1/A dadda_fa_2_79_1/B dadda_fa_2_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/CIN dadda_fa_3_79_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_56_0 dadda_fa_5_56_0/A dadda_fa_5_56_0/B dadda_fa_5_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/A dadda_fa_6_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_55_8 dadda_fa_1_55_8/A dadda_fa_1_55_8/B dadda_fa_1_55_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_56_3/A dadda_fa_3_55_0/A sky130_fd_sc_hd__fa_2
XFILLER_23_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_102_0 _694__914/HI U$$2738/X U$$2871/X VGND VGND VPWR VPWR dadda_fa_3_103_2/A
+ dadda_fa_3_102_3/A sky130_fd_sc_hd__fa_1
XFILLER_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1090 U$$1090/A _631_/Q VGND VGND VPWR VPWR U$$1090/X sky130_fd_sc_hd__xor2_1
XFILLER_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_81_1 U$$1632/X U$$1765/X U$$1898/X VGND VGND VPWR VPWR dadda_fa_2_82_1/B
+ dadda_fa_2_81_4/A sky130_fd_sc_hd__fa_1
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_74_0 U$$1751/X U$$1884/X U$$2017/X VGND VGND VPWR VPWR dadda_fa_2_75_0/B
+ dadda_fa_2_74_3/B sky130_fd_sc_hd__fa_2
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3409 U$$3409/A _665_/Q VGND VGND VPWR VPWR U$$3409/X sky130_fd_sc_hd__xor2_1
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2708 U$$2708/A _655_/Q VGND VGND VPWR VPWR U$$2708/X sky130_fd_sc_hd__xor2_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2719 _606_/Q U$$2607/X _607_/Q U$$2608/X VGND VGND VPWR VPWR U$$2720/A sky130_fd_sc_hd__a22o_1
XFILLER_74_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _611_/CLK _412_/D VGND VGND VPWR VPWR _412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _469_/CLK _343_/D VGND VGND VPWR VPWR _343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_274_ _280_/CLK _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_771__823 VGND VGND VPWR VPWR _771__823/HI U$$4389/B1 sky130_fd_sc_hd__conb_1
XFILLER_127_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_96_1 dadda_fa_3_96_1/A dadda_fa_3_96_1/B dadda_fa_3_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/CIN dadda_fa_4_96_2/A sky130_fd_sc_hd__fa_1
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_73_0 dadda_fa_6_73_0/A dadda_fa_6_73_0/B dadda_fa_6_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_74_0/B dadda_fa_7_73_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_6_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_89_0 dadda_fa_3_89_0/A dadda_fa_3_89_0/B dadda_fa_3_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/B dadda_fa_4_89_1/CIN sky130_fd_sc_hd__fa_1
X_812__864 VGND VGND VPWR VPWR _812__864/HI U$$4469/B sky130_fd_sc_hd__conb_1
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3910 _585_/Q U$$3840/X _586_/Q U$$3841/X VGND VGND VPWR VPWR U$$3911/A sky130_fd_sc_hd__a22o_1
XU$$3921 U$$3921/A _673_/Q VGND VGND VPWR VPWR U$$3921/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_118_0 _701__921/HI U$$3834/X U$$3967/X VGND VGND VPWR VPWR dadda_fa_5_119_0/B
+ dadda_fa_5_118_1/A sky130_fd_sc_hd__fa_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3932 _596_/Q U$$3970/A2 U$$98/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3933/A sky130_fd_sc_hd__a22o_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3943 U$$3943/A U$$3969/B VGND VGND VPWR VPWR U$$3943/X sky130_fd_sc_hd__xor2_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3954 U$$4502/A1 U$$3970/A2 U$$4504/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3955/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3965 U$$3965/A U$$3969/B VGND VGND VPWR VPWR U$$3965/X sky130_fd_sc_hd__xor2_2
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_5_5_0 U$$17/X U$$150/X VGND VGND VPWR VPWR dadda_fa_6_6_0/B dadda_fa_7_5_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_91_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3976 U$$4058/B U$$3976/B VGND VGND VPWR VPWR U$$3976/X sky130_fd_sc_hd__and2_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3987 U$$14/A1 U$$3977/X _556_/Q U$$3978/X VGND VGND VPWR VPWR U$$3988/A sky130_fd_sc_hd__a22o_1
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3998 U$$3998/A U$$4044/B VGND VGND VPWR VPWR U$$3998/X sky130_fd_sc_hd__xor2_1
XU$$170 U$$170/A U$$262/B VGND VGND VPWR VPWR U$$170/X sky130_fd_sc_hd__xor2_1
XFILLER_73_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$181 _570_/Q U$$141/X U$$46/A1 U$$142/X VGND VGND VPWR VPWR U$$182/A sky130_fd_sc_hd__a22o_1
XU$$192 U$$192/A U$$262/B VGND VGND VPWR VPWR U$$192/X sky130_fd_sc_hd__xor2_1
XFILLER_33_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_91_0 U$$3115/X U$$3248/X U$$3381/X VGND VGND VPWR VPWR dadda_fa_3_92_0/B
+ dadda_fa_3_91_2/B sky130_fd_sc_hd__fa_2
XFILLER_160_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput267 _277_/Q VGND VGND VPWR VPWR o[109] sky130_fd_sc_hd__buf_2
XFILLER_114_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput278 _287_/Q VGND VGND VPWR VPWR o[119] sky130_fd_sc_hd__buf_2
Xoutput289 _181_/Q VGND VGND VPWR VPWR o[13] sky130_fd_sc_hd__buf_2
XFILLER_142_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_47_6 U$$2495/X U$$2628/X VGND VGND VPWR VPWR dadda_fa_2_48_3/B dadda_fa_3_47_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_60_6 input213/X dadda_fa_1_60_6/B dadda_fa_1_60_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_61_2/B dadda_fa_2_60_5/B sky130_fd_sc_hd__fa_2
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_53_5 U$$2374/X U$$2507/X U$$2640/X VGND VGND VPWR VPWR dadda_fa_2_54_2/A
+ dadda_fa_2_53_5/A sky130_fd_sc_hd__fa_1
XFILLER_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_46_4 U$$1695/X U$$1828/X U$$1961/X VGND VGND VPWR VPWR dadda_fa_2_47_3/A
+ dadda_fa_2_46_5/B sky130_fd_sc_hd__fa_1
XFILLER_71_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_16_2 dadda_fa_4_16_2/A dadda_fa_4_16_2/B dadda_ha_3_16_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_17_0/CIN dadda_fa_5_16_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_755__807 VGND VGND VPWR VPWR _755__807/HI U$$3833/B1 sky130_fd_sc_hd__conb_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_90_0 dadda_fa_7_90_0/A dadda_fa_7_90_0/B dadda_fa_7_90_0/CIN VGND VGND
+ VPWR VPWR _515_/D _386_/D sky130_fd_sc_hd__fa_1
XFILLER_165_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3206 U$$3206/A U$$3244/B VGND VGND VPWR VPWR U$$3206/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3217 U$$3489/B1 U$$3241/A2 U$$3217/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3218/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3228 U$$3228/A U$$3244/B VGND VGND VPWR VPWR U$$3228/X sky130_fd_sc_hd__xor2_1
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3239 U$$771/B1 U$$3241/A2 U$$912/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3240/A sky130_fd_sc_hd__a22o_1
XFILLER_98_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2505 U$$2505/A U$$2533/B VGND VGND VPWR VPWR U$$2505/X sky130_fd_sc_hd__xor2_1
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2516 _573_/Q U$$2584/A2 U$$50/B1 U$$2584/B2 VGND VGND VPWR VPWR U$$2517/A sky130_fd_sc_hd__a22o_1
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2527 U$$2527/A U$$2585/B VGND VGND VPWR VPWR U$$2527/X sky130_fd_sc_hd__xor2_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2538 U$$892/B1 U$$2584/A2 U$$74/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2539/A sky130_fd_sc_hd__a22o_1
XU$$1804 U$$1804/A U$$1856/B VGND VGND VPWR VPWR U$$1804/X sky130_fd_sc_hd__xor2_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2549 U$$2549/A U$$2603/A VGND VGND VPWR VPWR U$$2549/X sky130_fd_sc_hd__xor2_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1815 U$$3457/B1 U$$1867/A2 U$$36/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1816/A sky130_fd_sc_hd__a22o_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1826 U$$1826/A U$$1872/B VGND VGND VPWR VPWR U$$1826/X sky130_fd_sc_hd__xor2_1
XU$$1837 U$$878/A1 U$$1903/A2 U$$880/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1838/A sky130_fd_sc_hd__a22o_1
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1848 U$$1848/A U$$1856/B VGND VGND VPWR VPWR U$$1848/X sky130_fd_sc_hd__xor2_1
XFILLER_42_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1859 U$$76/B1 U$$1897/A2 U$$902/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1860/A sky130_fd_sc_hd__a22o_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_326_ _339_/CLK _326_/D VGND VGND VPWR VPWR _326_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_257_ _267_/CLK _257_/D VGND VGND VPWR VPWR _257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_188_ _329_/CLK _188_/D VGND VGND VPWR VPWR _188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_70_5 dadda_fa_2_70_5/A dadda_fa_2_70_5/B dadda_fa_2_70_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_2/A dadda_fa_4_70_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_63_4 dadda_fa_2_63_4/A dadda_fa_2_63_4/B dadda_fa_2_63_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/CIN dadda_fa_3_63_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater704 U$$4303/A1 VGND VGND VPWR VPWR U$$878/A1 sky130_fd_sc_hd__buf_12
Xrepeater715 U$$4156/B1 VGND VGND VPWR VPWR U$$48/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater726 _568_/Q VGND VGND VPWR VPWR U$$4424/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_56_3 dadda_fa_2_56_3/A dadda_fa_2_56_3/B dadda_fa_2_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/B dadda_fa_3_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_42_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater737 U$$28/A1 VGND VGND VPWR VPWR U$$987/A1 sky130_fd_sc_hd__buf_12
XFILLER_111_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4430 _571_/Q U$$4388/X _572_/Q U$$4389/X VGND VGND VPWR VPWR U$$4431/A sky130_fd_sc_hd__a22o_1
Xrepeater748 U$$4265/A1 VGND VGND VPWR VPWR U$$18/A1 sky130_fd_sc_hd__buf_12
XU$$4441 U$$4441/A U$$4441/B VGND VGND VPWR VPWR U$$4441/X sky130_fd_sc_hd__xor2_4
Xrepeater759 _553_/Q VGND VGND VPWR VPWR U$$969/A1 sky130_fd_sc_hd__buf_12
XU$$4452 _582_/Q U$$4388/X U$$70/A1 U$$4389/X VGND VGND VPWR VPWR U$$4453/A sky130_fd_sc_hd__a22o_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_49_2 dadda_fa_2_49_2/A dadda_fa_2_49_2/B dadda_fa_2_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/A dadda_fa_3_49_3/A sky130_fd_sc_hd__fa_1
XU$$4463 U$$4463/A U$$4463/B VGND VGND VPWR VPWR U$$4463/X sky130_fd_sc_hd__xor2_2
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4474 U$$90/A1 U$$4388/X U$$4476/A1 U$$4389/X VGND VGND VPWR VPWR U$$4475/A sky130_fd_sc_hd__a22o_1
XU$$3740 U$$3740/A U$$3756/B VGND VGND VPWR VPWR U$$3740/X sky130_fd_sc_hd__xor2_1
XU$$4485 U$$4485/A U$$4485/B VGND VGND VPWR VPWR U$$4485/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_26_1 dadda_fa_5_26_1/A dadda_fa_5_26_1/B dadda_fa_5_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/B dadda_fa_7_26_0/A sky130_fd_sc_hd__fa_1
XFILLER_93_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3751 _574_/Q U$$3795/A2 _575_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3752/A sky130_fd_sc_hd__a22o_1
XU$$4496 U$$4496/A1 U$$4388/X U$$936/A1 U$$4389/X VGND VGND VPWR VPWR U$$4497/A sky130_fd_sc_hd__a22o_1
XFILLER_65_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3762 U$$3762/A U$$3794/B VGND VGND VPWR VPWR U$$3762/X sky130_fd_sc_hd__xor2_1
XFILLER_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3773 _585_/Q U$$3795/A2 _586_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3774/A sky130_fd_sc_hd__a22o_1
XFILLER_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_19_0 dadda_fa_5_19_0/A dadda_fa_5_19_0/B dadda_fa_5_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/A dadda_fa_6_19_0/CIN sky130_fd_sc_hd__fa_1
XU$$3784 U$$3784/A U$$3784/B VGND VGND VPWR VPWR U$$3784/X sky130_fd_sc_hd__xor2_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3795 U$$96/A1 U$$3795/A2 _597_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3796/A sky130_fd_sc_hd__a22o_1
XFILLER_166_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_100_1 dadda_fa_5_100_1/A dadda_fa_5_100_1/B dadda_fa_5_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/B dadda_fa_7_100_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_122_0 _708__928/HI U$$4108/X VGND VGND VPWR VPWR dadda_fa_5_123_1/CIN
+ dadda_ha_4_122_0/SUM sky130_fd_sc_hd__ha_1
XFILLER_86_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_1_38_2 U$$881/X U$$1014/X VGND VGND VPWR VPWR dadda_fa_2_39_5/A dadda_fa_3_38_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_134_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_51_2 U$$907/X U$$1040/X U$$1173/X VGND VGND VPWR VPWR dadda_fa_2_52_1/A
+ dadda_fa_2_51_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$906 U$$84/A1 U$$928/A2 U$$908/A1 U$$928/B2 VGND VGND VPWR VPWR U$$907/A sky130_fd_sc_hd__a22o_1
XFILLER_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$917 U$$917/A U$$943/B VGND VGND VPWR VPWR U$$917/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_1 U$$494/X U$$627/X U$$760/X VGND VGND VPWR VPWR dadda_fa_2_45_2/CIN
+ dadda_fa_2_44_4/CIN sky130_fd_sc_hd__fa_2
XU$$928 U$$928/A1 U$$928/A2 U$$928/B1 U$$928/B2 VGND VGND VPWR VPWR U$$929/A sky130_fd_sc_hd__a22o_1
XFILLER_56_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$939 U$$939/A _629_/Q VGND VGND VPWR VPWR U$$939/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_21_0 input170/X dadda_fa_4_21_0/B dadda_fa_4_21_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_22_0/A dadda_fa_5_21_1/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_37_0 U$$81/X U$$214/X U$$347/X VGND VGND VPWR VPWR dadda_fa_2_38_4/CIN
+ dadda_fa_2_37_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_73_3 dadda_fa_3_73_3/A dadda_fa_3_73_3/B dadda_fa_3_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/B dadda_fa_4_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_66_2 dadda_fa_3_66_2/A dadda_fa_3_66_2/B dadda_fa_3_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/A dadda_fa_4_66_2/B sky130_fd_sc_hd__fa_1
XFILLER_132_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_59_1 dadda_fa_3_59_1/A dadda_fa_3_59_1/B dadda_fa_3_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/CIN dadda_fa_4_59_2/A sky130_fd_sc_hd__fa_1
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_36_0 dadda_fa_6_36_0/A dadda_fa_6_36_0/B dadda_fa_6_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_37_0/B dadda_fa_7_36_0/CIN sky130_fd_sc_hd__fa_2
XU$$3003 _611_/Q U$$2881/X _612_/Q U$$2882/X VGND VGND VPWR VPWR U$$3004/A sky130_fd_sc_hd__a22o_1
XU$$3014 _659_/Q VGND VGND VPWR VPWR U$$3014/Y sky130_fd_sc_hd__inv_1
XU$$3025 U$$3025/A U$$3085/B VGND VGND VPWR VPWR U$$3025/X sky130_fd_sc_hd__xor2_1
XU$$3036 U$$979/B1 U$$3090/A2 U$$4271/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3037/A
+ sky130_fd_sc_hd__a22o_1
XU$$2302 _603_/Q U$$2326/A2 _604_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2303/A sky130_fd_sc_hd__a22o_1
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3047 U$$3047/A U$$3085/B VGND VGND VPWR VPWR U$$3047/X sky130_fd_sc_hd__xor2_1
XU$$2313 U$$2313/A _649_/Q VGND VGND VPWR VPWR U$$2313/X sky130_fd_sc_hd__xor2_1
XU$$3058 U$$4291/A1 U$$3146/A2 U$$868/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3059/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2324 U$$4379/A1 U$$2196/X U$$819/A1 U$$2197/X VGND VGND VPWR VPWR U$$2325/A sky130_fd_sc_hd__a22o_1
XFILLER_74_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3069 U$$3069/A U$$3085/B VGND VGND VPWR VPWR U$$3069/X sky130_fd_sc_hd__xor2_1
XU$$2335 U$$2335/A1 U$$2333/X U$$8/A1 U$$2334/X VGND VGND VPWR VPWR U$$2336/A sky130_fd_sc_hd__a22o_1
XU$$1601 U$$94/A1 U$$1511/X U$$94/B1 U$$1512/X VGND VGND VPWR VPWR U$$1602/A sky130_fd_sc_hd__a22o_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2346 U$$2346/A U$$2432/B VGND VGND VPWR VPWR U$$2346/X sky130_fd_sc_hd__xor2_1
XU$$2357 U$$28/A1 U$$2421/A2 U$$30/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2358/A sky130_fd_sc_hd__a22o_1
XFILLER_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1612 U$$1612/A _639_/Q VGND VGND VPWR VPWR U$$1612/X sky130_fd_sc_hd__xor2_1
XU$$1623 _606_/Q U$$1641/A2 _607_/Q U$$1641/B2 VGND VGND VPWR VPWR U$$1624/A sky130_fd_sc_hd__a22o_1
XU$$2368 U$$2368/A U$$2436/B VGND VGND VPWR VPWR U$$2368/X sky130_fd_sc_hd__xor2_1
XU$$2379 _573_/Q U$$2421/A2 U$$2790/B1 U$$2421/B2 VGND VGND VPWR VPWR U$$2380/A sky130_fd_sc_hd__a22o_1
XU$$1634 U$$1634/A _639_/Q VGND VGND VPWR VPWR U$$1634/X sky130_fd_sc_hd__xor2_1
XU$$1645 _640_/Q VGND VGND VPWR VPWR U$$1647/B sky130_fd_sc_hd__inv_1
XFILLER_43_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1656 U$$12/A1 U$$1734/A2 U$$14/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1657/A sky130_fd_sc_hd__a22o_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1667 U$$1667/A U$$1727/B VGND VGND VPWR VPWR U$$1667/X sky130_fd_sc_hd__xor2_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1678 U$$3457/B1 U$$1734/A2 U$$36/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1679/A sky130_fd_sc_hd__a22o_1
XFILLER_187_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1689 U$$1689/A U$$1727/B VGND VGND VPWR VPWR U$$1689/X sky130_fd_sc_hd__xor2_1
XFILLER_129_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_309_ _463_/CLK _309_/D VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_818__870 VGND VGND VPWR VPWR _818__870/HI U$$4481/B sky130_fd_sc_hd__conb_1
Xdadda_fa_7_109_0 dadda_fa_7_109_0/A dadda_fa_7_109_0/B dadda_fa_7_109_0/CIN VGND
+ VGND VPWR VPWR _534_/D _405_/D sky130_fd_sc_hd__fa_2
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_61_1 dadda_fa_2_61_1/A dadda_fa_2_61_1/B dadda_fa_2_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/CIN dadda_fa_3_61_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater501 U$$1786/X VGND VGND VPWR VPWR U$$1897/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$308 final_adder.U$$308/A final_adder.U$$308/B VGND VGND VPWR VPWR
+ final_adder.U$$346/B sky130_fd_sc_hd__and2_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater512 U$$1238/X VGND VGND VPWR VPWR U$$1367/B2 sky130_fd_sc_hd__buf_12
XFILLER_111_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater523 _673_/Q VGND VGND VPWR VPWR U$$3929/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_54_0 dadda_fa_2_54_0/A dadda_fa_2_54_0/B dadda_fa_2_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/B dadda_fa_3_54_2/B sky130_fd_sc_hd__fa_2
Xrepeater534 U$$3536/B VGND VGND VPWR VPWR U$$3496/B sky130_fd_sc_hd__buf_12
Xrepeater545 _661_/Q VGND VGND VPWR VPWR U$$3137/B sky130_fd_sc_hd__buf_12
XFILLER_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater556 _653_/Q VGND VGND VPWR VPWR U$$2585/B sky130_fd_sc_hd__buf_12
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater567 U$$2023/B VGND VGND VPWR VPWR U$$1991/B sky130_fd_sc_hd__buf_12
XU$$4260 U$$4260/A U$$4384/A VGND VGND VPWR VPWR U$$4260/X sky130_fd_sc_hd__xor2_1
Xrepeater578 U$$1614/B VGND VGND VPWR VPWR U$$1580/B sky130_fd_sc_hd__buf_12
XFILLER_26_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4271 U$$4271/A1 U$$4381/A2 _561_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4272/A sky130_fd_sc_hd__a22o_1
Xrepeater589 _633_/Q VGND VGND VPWR VPWR U$$1232/A sky130_fd_sc_hd__buf_12
XU$$4282 U$$4282/A U$$4384/A VGND VGND VPWR VPWR U$$4282/X sky130_fd_sc_hd__xor2_1
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4293 _571_/Q U$$4377/A2 _572_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4294/A sky130_fd_sc_hd__a22o_1
XFILLER_77_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3570 U$$4255/A1 U$$3624/A2 U$$969/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3571/A
+ sky130_fd_sc_hd__a22o_1
XU$$3581 U$$3581/A U$$3625/B VGND VGND VPWR VPWR U$$3581/X sky130_fd_sc_hd__xor2_1
XU$$3592 _563_/Q U$$3678/A2 U$$32/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3593/A sky130_fd_sc_hd__a22o_1
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_8_0 U$$289/X U$$422/X U$$555/X VGND VGND VPWR VPWR dadda_fa_6_9_0/A dadda_fa_6_8_0/CIN
+ sky130_fd_sc_hd__fa_2
XU$$2880 _659_/Q U$$2880/B VGND VGND VPWR VPWR U$$2880/X sky130_fd_sc_hd__and2_1
XFILLER_80_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2891 U$$14/A1 U$$3009/A2 U$$14/B1 U$$3009/B2 VGND VGND VPWR VPWR U$$2892/A sky130_fd_sc_hd__a22o_1
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_83_2 dadda_fa_4_83_2/A dadda_fa_4_83_2/B dadda_fa_4_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/CIN dadda_fa_5_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_76_1 dadda_fa_4_76_1/A dadda_fa_4_76_1/B dadda_fa_4_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/B dadda_fa_5_76_1/B sky130_fd_sc_hd__fa_1
XFILLER_136_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_53_0 dadda_fa_7_53_0/A dadda_fa_7_53_0/B dadda_fa_7_53_0/CIN VGND VGND
+ VPWR VPWR _478_/D _349_/D sky130_fd_sc_hd__fa_2
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_69_0 dadda_fa_4_69_0/A dadda_fa_4_69_0/B dadda_fa_4_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/A dadda_fa_5_69_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_660_ _667_/CLK _660_/D VGND VGND VPWR VPWR _660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$703 U$$18/A1 U$$817/A2 U$$842/A1 U$$785/B2 VGND VGND VPWR VPWR U$$704/A sky130_fd_sc_hd__a22o_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$714 U$$714/A U$$778/B VGND VGND VPWR VPWR U$$714/X sky130_fd_sc_hd__xor2_1
XFILLER_112_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$725 U$$40/A1 U$$817/A2 _569_/Q U$$785/B2 VGND VGND VPWR VPWR U$$726/A sky130_fd_sc_hd__a22o_1
X_591_ _595_/CLK _591_/D VGND VGND VPWR VPWR _591_/Q sky130_fd_sc_hd__dfxtp_4
XU$$736 U$$736/A U$$784/B VGND VGND VPWR VPWR U$$736/X sky130_fd_sc_hd__xor2_1
XFILLER_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$747 U$$62/A1 U$$689/X U$$64/A1 U$$817/B2 VGND VGND VPWR VPWR U$$748/A sky130_fd_sc_hd__a22o_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$758 U$$758/A U$$778/B VGND VGND VPWR VPWR U$$758/X sky130_fd_sc_hd__xor2_1
XU$$769 U$$84/A1 U$$785/A2 U$$86/A1 U$$785/B2 VGND VGND VPWR VPWR U$$770/A sky130_fd_sc_hd__a22o_1
XFILLER_32_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_71_0 dadda_fa_3_71_0/A dadda_fa_3_71_0/B dadda_fa_3_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/B dadda_fa_4_71_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2110 U$$2110/A U$$2118/B VGND VGND VPWR VPWR U$$2110/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_100_0 dadda_fa_4_100_0/A dadda_fa_4_100_0/B dadda_fa_4_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/A dadda_fa_5_100_1/A sky130_fd_sc_hd__fa_1
XU$$2121 U$$3489/B1 U$$2161/A2 U$$3217/B1 U$$2161/B2 VGND VGND VPWR VPWR U$$2122/A
+ sky130_fd_sc_hd__a22o_1
XU$$2132 U$$2132/A U$$2186/B VGND VGND VPWR VPWR U$$2132/X sky130_fd_sc_hd__xor2_1
XU$$2143 U$$4335/A1 U$$2161/A2 _593_/Q U$$2161/B2 VGND VGND VPWR VPWR U$$2144/A sky130_fd_sc_hd__a22o_1
XU$$2154 U$$2154/A U$$2192/A VGND VGND VPWR VPWR U$$2154/X sky130_fd_sc_hd__xor2_1
XU$$1420 U$$735/A1 U$$1474/A2 U$$52/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1421/A sky130_fd_sc_hd__a22o_1
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2165 _603_/Q U$$2189/A2 U$$4496/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2166/A sky130_fd_sc_hd__a22o_1
XU$$2176 U$$2176/A U$$2192/A VGND VGND VPWR VPWR U$$2176/X sky130_fd_sc_hd__xor2_1
XU$$1431 U$$1431/A U$$1461/B VGND VGND VPWR VPWR U$$1431/X sky130_fd_sc_hd__xor2_1
XU$$1442 U$$892/B1 U$$1472/A2 U$$74/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1443/A sky130_fd_sc_hd__a22o_1
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2187 _614_/Q U$$2189/A2 _615_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2188/A sky130_fd_sc_hd__a22o_1
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2198 U$$2198/A1 U$$2196/X U$$8/A1 U$$2197/X VGND VGND VPWR VPWR U$$2199/A sky130_fd_sc_hd__a22o_1
XU$$1453 U$$1453/A U$$1505/B VGND VGND VPWR VPWR U$$1453/X sky130_fd_sc_hd__xor2_1
XU$$1464 U$$94/A1 U$$1474/A2 U$$94/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1465/A sky130_fd_sc_hd__a22o_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1475 U$$1475/A U$$1479/B VGND VGND VPWR VPWR U$$1475/X sky130_fd_sc_hd__xor2_1
XFILLER_176_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1486 U$$938/A1 U$$1374/X _607_/Q U$$1375/X VGND VGND VPWR VPWR U$$1487/A sky130_fd_sc_hd__a22o_1
XFILLER_187_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1497 U$$1497/A _637_/Q VGND VGND VPWR VPWR U$$1497/X sky130_fd_sc_hd__xor2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_93_1 dadda_fa_5_93_1/A dadda_fa_5_93_1/B dadda_fa_5_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/B dadda_fa_7_93_0/A sky130_fd_sc_hd__fa_2
XFILLER_191_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_86_0 dadda_fa_5_86_0/A dadda_fa_5_86_0/B dadda_fa_5_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/A dadda_fa_6_86_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_7 U$$4020/X U$$4153/X U$$4286/X VGND VGND VPWR VPWR dadda_fa_2_79_2/CIN
+ dadda_fa_2_78_5/CIN sky130_fd_sc_hd__fa_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$105 _529_/Q _401_/Q VGND VGND VPWR VPWR final_adder.U$$233/B1 final_adder.U$$727/A
+ sky130_fd_sc_hd__ha_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$116 _540_/Q _412_/Q VGND VGND VPWR VPWR final_adder.U$$611/B1 final_adder.U$$738/A
+ sky130_fd_sc_hd__ha_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$127 _551_/Q _423_/Q VGND VGND VPWR VPWR final_adder.U$$127/COUT final_adder.U$$749/A
+ sky130_fd_sc_hd__ha_4
XFILLER_170_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$138 final_adder.U$$633/A final_adder.U$$632/A VGND VGND VPWR VPWR
+ final_adder.U$$260/A sky130_fd_sc_hd__and2_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$149 final_adder.U$$643/A final_adder.U$$515/B1 final_adder.U$$149/B1
+ VGND VGND VPWR VPWR final_adder.U$$149/X sky130_fd_sc_hd__a21o_1
XFILLER_38_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater386 U$$963/X VGND VGND VPWR VPWR U$$1093/A2 sky130_fd_sc_hd__buf_12
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater397 U$$4114/X VGND VGND VPWR VPWR U$$4244/A2 sky130_fd_sc_hd__buf_12
XU$$4090 U$$4090/A U$$4109/A VGND VGND VPWR VPWR U$$4090/X sky130_fd_sc_hd__xor2_1
XFILLER_54_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_102_2 dadda_fa_3_102_2/A dadda_fa_3_102_2/B dadda_fa_3_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/A dadda_fa_4_102_2/B sky130_fd_sc_hd__fa_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput101 b[42] VGND VGND VPWR VPWR _594_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput112 b[52] VGND VGND VPWR VPWR _604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput123 b[62] VGND VGND VPWR VPWR _614_/D sky130_fd_sc_hd__clkbuf_4
Xinput134 c[104] VGND VGND VPWR VPWR input134/X sky130_fd_sc_hd__buf_2
Xinput145 c[114] VGND VGND VPWR VPWR input145/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_66_5 U$$2134/X U$$2267/X U$$2400/X VGND VGND VPWR VPWR dadda_fa_1_67_7/A
+ dadda_fa_2_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput156 c[124] VGND VGND VPWR VPWR input156/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 c[19] VGND VGND VPWR VPWR input167/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_6_116_0 dadda_fa_6_116_0/A dadda_fa_6_116_0/B dadda_fa_6_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_117_0/B dadda_fa_7_116_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput178 c[29] VGND VGND VPWR VPWR input178/X sky130_fd_sc_hd__clkbuf_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 c[39] VGND VGND VPWR VPWR input189/X sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$650 final_adder.U$$650/A final_adder.U$$650/B VGND VGND VPWR VPWR
+ _196_/D sky130_fd_sc_hd__xor2_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$661 final_adder.U$$661/A final_adder.U$$661/B VGND VGND VPWR VPWR
+ _207_/D sky130_fd_sc_hd__xor2_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$500 U$$500/A _623_/Q VGND VGND VPWR VPWR U$$500/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$672 final_adder.U$$672/A final_adder.U$$672/B VGND VGND VPWR VPWR
+ _218_/D sky130_fd_sc_hd__xor2_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_643_ _647_/CLK _643_/D VGND VGND VPWR VPWR _643_/Q sky130_fd_sc_hd__dfxtp_4
XU$$511 U$$785/A1 U$$545/A2 U$$924/A1 U$$416/X VGND VGND VPWR VPWR U$$512/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_36_3 dadda_fa_3_36_3/A dadda_fa_3_36_3/B dadda_fa_3_36_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/B dadda_fa_4_36_2/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$683 final_adder.U$$683/A final_adder.U$$683/B VGND VGND VPWR VPWR
+ _229_/D sky130_fd_sc_hd__xor2_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$522 U$$522/A U$$547/A VGND VGND VPWR VPWR U$$522/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$694 final_adder.U$$694/A final_adder.U$$694/B VGND VGND VPWR VPWR
+ _240_/D sky130_fd_sc_hd__xor2_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$533 U$$944/A1 U$$415/X U$$946/A1 U$$416/X VGND VGND VPWR VPWR U$$534/A sky130_fd_sc_hd__a22o_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$544 U$$544/A U$$547/A VGND VGND VPWR VPWR U$$544/X sky130_fd_sc_hd__xor2_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$555 U$$555/A U$$623/B VGND VGND VPWR VPWR U$$555/X sky130_fd_sc_hd__xor2_1
XFILLER_44_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_29_2 dadda_fa_3_29_2/A dadda_fa_3_29_2/B dadda_fa_3_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/A dadda_fa_4_29_2/B sky130_fd_sc_hd__fa_2
XU$$566 U$$18/A1 U$$626/A2 U$$20/A1 U$$553/X VGND VGND VPWR VPWR U$$567/A sky130_fd_sc_hd__a22o_1
XFILLER_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_574_ _679_/CLK _574_/D VGND VGND VPWR VPWR _574_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$577 U$$577/A U$$623/B VGND VGND VPWR VPWR U$$577/X sky130_fd_sc_hd__xor2_1
XU$$588 U$$40/A1 U$$626/A2 _569_/Q U$$553/X VGND VGND VPWR VPWR U$$589/A sky130_fd_sc_hd__a22o_1
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$599 U$$599/A U$$623/B VGND VGND VPWR VPWR U$$599/X sky130_fd_sc_hd__xor2_1
XFILLER_112_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_31_2 U$$867/X U$$1000/X U$$1133/X VGND VGND VPWR VPWR dadda_fa_3_32_1/B
+ dadda_fa_3_31_3/B sky130_fd_sc_hd__fa_1
XFILLER_51_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1250 U$$1250/A U$$1336/B VGND VGND VPWR VPWR U$$1250/X sky130_fd_sc_hd__xor2_1
XFILLER_189_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1261 U$$28/A1 U$$1237/X U$$28/B1 U$$1238/X VGND VGND VPWR VPWR U$$1262/A sky130_fd_sc_hd__a22o_1
XU$$1272 U$$1272/A U$$1342/B VGND VGND VPWR VPWR U$$1272/X sky130_fd_sc_hd__xor2_1
XFILLER_188_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1283 U$$50/A1 U$$1341/A2 U$$50/B1 U$$1341/B2 VGND VGND VPWR VPWR U$$1284/A sky130_fd_sc_hd__a22o_1
XU$$1294 U$$1294/A U$$1342/B VGND VGND VPWR VPWR U$$1294/X sky130_fd_sc_hd__xor2_1
XFILLER_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_5 U$$3365/X U$$3498/X U$$3631/X VGND VGND VPWR VPWR dadda_fa_2_84_3/B
+ dadda_fa_2_83_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_116_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_76_4 U$$3085/X U$$3218/X U$$3351/X VGND VGND VPWR VPWR dadda_fa_2_77_1/CIN
+ dadda_fa_2_76_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_3 U$$3603/X U$$3736/X U$$3869/X VGND VGND VPWR VPWR dadda_fa_2_70_1/B
+ dadda_fa_2_69_4/B sky130_fd_sc_hd__fa_1
XFILLER_140_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_46_2 dadda_fa_4_46_2/A dadda_fa_4_46_2/B dadda_fa_4_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/CIN dadda_fa_5_46_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_1 dadda_fa_4_39_1/A dadda_fa_4_39_1/B dadda_fa_4_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/B dadda_fa_5_39_1/B sky130_fd_sc_hd__fa_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_16_0 dadda_fa_7_16_0/A dadda_fa_7_16_0/B dadda_fa_7_16_0/CIN VGND VGND
+ VPWR VPWR _441_/D _312_/D sky130_fd_sc_hd__fa_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_723__775 VGND VGND VPWR VPWR _723__775/HI U$$1778/B1 sky130_fd_sc_hd__conb_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ _612_/CLK _290_/D VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_0_58_3 U$$1320/X U$$1453/X VGND VGND VPWR VPWR dadda_fa_1_59_7/CIN dadda_fa_2_58_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_71_3 U$$1745/X U$$1878/X U$$2011/X VGND VGND VPWR VPWR dadda_fa_1_72_7/CIN
+ dadda_fa_2_71_0/A sky130_fd_sc_hd__fa_2
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_64_2 U$$933/X U$$1066/X U$$1199/X VGND VGND VPWR VPWR dadda_fa_1_65_6/A
+ dadda_fa_1_64_8/A sky130_fd_sc_hd__fa_1
XFILLER_114_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_41_1 dadda_fa_3_41_1/A dadda_fa_3_41_1/B dadda_fa_3_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/CIN dadda_fa_4_41_2/A sky130_fd_sc_hd__fa_2
XFILLER_188_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_57_1 U$$520/X U$$653/X U$$786/X VGND VGND VPWR VPWR dadda_fa_1_58_7/B
+ dadda_fa_1_57_8/CIN sky130_fd_sc_hd__fa_2
XFILLER_188_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_34_0 dadda_fa_3_34_0/A dadda_fa_3_34_0/B dadda_fa_3_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/B dadda_fa_4_34_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$491 final_adder.U$$314/B final_adder.U$$738/B final_adder.U$$245/X
+ VGND VGND VPWR VPWR final_adder.U$$740/B sky130_fd_sc_hd__a21o_1
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$330 U$$56/A1 U$$278/X U$$58/A1 U$$279/X VGND VGND VPWR VPWR U$$331/A sky130_fd_sc_hd__a22o_1
X_626_ _633_/CLK _626_/D VGND VGND VPWR VPWR _626_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$341 U$$341/A U$$357/B VGND VGND VPWR VPWR U$$341/X sky130_fd_sc_hd__xor2_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$352 U$$78/A1 U$$278/X U$$80/A1 U$$279/X VGND VGND VPWR VPWR U$$353/A sky130_fd_sc_hd__a22o_1
XFILLER_18_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$363 U$$363/A _621_/Q VGND VGND VPWR VPWR U$$363/X sky130_fd_sc_hd__xor2_1
XU$$374 U$$785/A1 U$$278/X U$$924/A1 U$$279/X VGND VGND VPWR VPWR U$$375/A sky130_fd_sc_hd__a22o_1
XU$$385 U$$385/A U$$391/B VGND VGND VPWR VPWR U$$385/X sky130_fd_sc_hd__xor2_1
XFILLER_72_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_557_ _649_/CLK _557_/D VGND VGND VPWR VPWR _557_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$396 U$$944/A1 U$$278/X U$$946/A1 U$$279/X VGND VGND VPWR VPWR U$$397/A sky130_fd_sc_hd__a22o_1
XFILLER_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_488_ _488_/CLK _488_/D VGND VGND VPWR VPWR _488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_93_4 U$$4449/X input249/X dadda_fa_2_93_4/CIN VGND VGND VPWR VPWR dadda_fa_3_94_1/CIN
+ dadda_fa_3_93_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_86_3 dadda_fa_2_86_3/A dadda_fa_2_86_3/B dadda_fa_2_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/B dadda_fa_3_86_3/B sky130_fd_sc_hd__fa_2
XFILLER_99_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_79_2 dadda_fa_2_79_2/A dadda_fa_2_79_2/B dadda_fa_2_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/A dadda_fa_3_79_3/A sky130_fd_sc_hd__fa_2
XFILLER_99_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_56_1 dadda_fa_5_56_1/A dadda_fa_5_56_1/B dadda_fa_5_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/B dadda_fa_7_56_0/A sky130_fd_sc_hd__fa_1
XFILLER_45_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_49_0 dadda_fa_5_49_0/A dadda_fa_5_49_0/B dadda_fa_5_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/A dadda_fa_6_49_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_23_0 U$$53/X U$$186/X VGND VGND VPWR VPWR dadda_fa_3_24_3/B dadda_fa_4_23_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_102_1 U$$3004/X U$$3137/X U$$3270/X VGND VGND VPWR VPWR dadda_fa_3_103_2/B
+ dadda_fa_3_102_3/B sky130_fd_sc_hd__fa_2
XFILLER_51_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1080 U$$1080/A _631_/Q VGND VGND VPWR VPWR U$$1080/X sky130_fd_sc_hd__xor2_1
XU$$1091 U$$952/B1 U$$963/X U$$819/A1 U$$964/X VGND VGND VPWR VPWR U$$1092/A sky130_fd_sc_hd__a22o_1
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_123_0 U$$4109/Y U$$4243/X U$$4376/X VGND VGND VPWR VPWR dadda_fa_6_124_0/A
+ dadda_fa_6_123_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_52_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk _369_/CLK VGND VGND VPWR VPWR _471_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_81_2 U$$2031/X U$$2164/X U$$2297/X VGND VGND VPWR VPWR dadda_fa_2_82_1/CIN
+ dadda_fa_2_81_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_74_1 U$$2150/X U$$2283/X U$$2416/X VGND VGND VPWR VPWR dadda_fa_2_75_0/CIN
+ dadda_fa_2_74_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_51_0 dadda_fa_4_51_0/A dadda_fa_4_51_0/B dadda_fa_4_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/A dadda_fa_5_51_1/A sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_97_clk _431_/CLK VGND VGND VPWR VPWR _432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_67_0 U$$2535/X U$$2668/X U$$2801/X VGND VGND VPWR VPWR dadda_fa_2_68_0/B
+ dadda_fa_2_67_3/B sky130_fd_sc_hd__fa_2
XFILLER_58_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2709 _601_/Q U$$2729/A2 U$$928/B1 U$$2729/B2 VGND VGND VPWR VPWR U$$2710/A sky130_fd_sc_hd__a22o_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _611_/CLK _411_/D VGND VGND VPWR VPWR _411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ _476_/CLK _342_/D VGND VGND VPWR VPWR _342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_273_ _280_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _329_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_96_2 dadda_fa_3_96_2/A dadda_fa_3_96_2/B dadda_fa_3_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/A dadda_fa_4_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_89_1 dadda_fa_3_89_1/A dadda_fa_3_89_1/B dadda_fa_3_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/CIN dadda_fa_4_89_2/A sky130_fd_sc_hd__fa_2
XFILLER_136_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_66_0 dadda_fa_6_66_0/A dadda_fa_6_66_0/B dadda_fa_6_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_67_0/B dadda_fa_7_66_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _649_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3900 U$$3900/A1 U$$3912/A2 _581_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3901/A sky130_fd_sc_hd__a22o_1
XU$$3911 U$$3911/A _673_/Q VGND VGND VPWR VPWR U$$3911/X sky130_fd_sc_hd__xor2_1
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_118_1 U$$4100/X U$$4233/X U$$4366/X VGND VGND VPWR VPWR dadda_fa_5_119_0/CIN
+ dadda_fa_5_118_1/B sky130_fd_sc_hd__fa_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3922 _591_/Q U$$3840/X U$$4335/A1 U$$3841/X VGND VGND VPWR VPWR U$$3923/A sky130_fd_sc_hd__a22o_1
XU$$3933 U$$3933/A _673_/Q VGND VGND VPWR VPWR U$$3933/X sky130_fd_sc_hd__xor2_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3944 U$$4492/A1 U$$3970/A2 U$$4494/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3945/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3955 U$$3955/A U$$3969/B VGND VGND VPWR VPWR U$$3955/X sky130_fd_sc_hd__xor2_1
XFILLER_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3966 _613_/Q U$$3970/A2 U$$4379/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3967/A sky130_fd_sc_hd__a22o_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3977 U$$3975/Y _674_/Q _673_/Q U$$3976/X U$$3973/Y VGND VGND VPWR VPWR U$$3977/X
+ sky130_fd_sc_hd__a32o_4
XU$$160 U$$160/A U$$274/A VGND VGND VPWR VPWR U$$160/X sky130_fd_sc_hd__xor2_1
XU$$3988 U$$3988/A U$$4058/B VGND VGND VPWR VPWR U$$3988/X sky130_fd_sc_hd__xor2_1
X_609_ _611_/CLK _609_/D VGND VGND VPWR VPWR _609_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3999 U$$4273/A1 U$$3977/X _562_/Q U$$3978/X VGND VGND VPWR VPWR U$$4000/A sky130_fd_sc_hd__a22o_1
XU$$171 U$$34/A1 U$$141/X U$$36/A1 U$$142/X VGND VGND VPWR VPWR U$$172/A sky130_fd_sc_hd__a22o_1
XFILLER_33_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$182 U$$182/A U$$242/B VGND VGND VPWR VPWR U$$182/X sky130_fd_sc_hd__xor2_1
XU$$193 U$$56/A1 U$$141/X U$$58/A1 U$$142/X VGND VGND VPWR VPWR U$$194/A sky130_fd_sc_hd__a22o_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_12_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _461_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_1 U$$3514/X U$$3647/X U$$3780/X VGND VGND VPWR VPWR dadda_fa_3_92_0/CIN
+ dadda_fa_3_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_84_0 U$$4032/X U$$4165/X U$$4298/X VGND VGND VPWR VPWR dadda_fa_3_85_0/B
+ dadda_fa_3_84_2/B sky130_fd_sc_hd__fa_2
XFILLER_160_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput257 _168_/Q VGND VGND VPWR VPWR o[0] sky130_fd_sc_hd__buf_2
XFILLER_82_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput268 _178_/Q VGND VGND VPWR VPWR o[10] sky130_fd_sc_hd__buf_2
Xoutput279 _179_/Q VGND VGND VPWR VPWR o[11] sky130_fd_sc_hd__buf_2
XFILLER_82_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_60_7 dadda_fa_1_60_7/A dadda_fa_1_60_7/B dadda_fa_1_60_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_2/CIN dadda_fa_2_60_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_53_6 U$$2773/X U$$2906/X U$$3039/X VGND VGND VPWR VPWR dadda_fa_2_54_2/B
+ dadda_fa_2_53_5/B sky130_fd_sc_hd__fa_1
XFILLER_95_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_46_5 U$$2094/X U$$2227/X U$$2360/X VGND VGND VPWR VPWR dadda_fa_2_47_3/B
+ dadda_fa_2_46_5/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_7_5_0 dadda_fa_7_5_0/A dadda_fa_7_5_0/B dadda_fa_7_5_0/CIN VGND VGND VPWR
+ VPWR _430_/D _301_/D sky130_fd_sc_hd__fa_1
XFILLER_64_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_794__846 VGND VGND VPWR VPWR _794__846/HI U$$4433/B sky130_fd_sc_hd__conb_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_83_0 dadda_fa_7_83_0/A dadda_fa_7_83_0/B dadda_fa_7_83_0/CIN VGND VGND
+ VPWR VPWR _508_/D _379_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_99_0 dadda_fa_4_99_0/A dadda_fa_4_99_0/B dadda_fa_4_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/A dadda_fa_5_99_1/A sky130_fd_sc_hd__fa_1
XFILLER_180_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_835__887 VGND VGND VPWR VPWR _835__887/HI U$$4515/B sky130_fd_sc_hd__conb_1
XFILLER_104_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3207 U$$4303/A1 U$$3243/A2 U$$4442/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3208/A
+ sky130_fd_sc_hd__a22o_1
X_729__781 VGND VGND VPWR VPWR _729__781/HI U$$2189/B1 sky130_fd_sc_hd__conb_1
XFILLER_98_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3218 U$$3218/A U$$3224/B VGND VGND VPWR VPWR U$$3218/X sky130_fd_sc_hd__xor2_1
XU$$3229 _587_/Q U$$3243/A2 U$$902/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3230/A sky130_fd_sc_hd__a22o_1
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2506 U$$3191/A1 U$$2534/A2 U$$4289/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2507/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2517 U$$2517/A U$$2585/B VGND VGND VPWR VPWR U$$2517/X sky130_fd_sc_hd__xor2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2528 U$$4446/A1 U$$2574/A2 U$$64/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2529/A sky130_fd_sc_hd__a22o_1
XFILLER_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2539 U$$2539/A U$$2585/B VGND VGND VPWR VPWR U$$2539/X sky130_fd_sc_hd__xor2_1
XU$$1805 U$$4271/A1 U$$1903/A2 U$$4273/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1806/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1816 U$$1816/A U$$1918/A VGND VGND VPWR VPWR U$$1816/X sky130_fd_sc_hd__xor2_1
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1827 U$$868/A1 U$$1897/A2 U$$48/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1828/A sky130_fd_sc_hd__a22o_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1838 U$$1838/A U$$1856/B VGND VGND VPWR VPWR U$$1838/X sky130_fd_sc_hd__xor2_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1849 U$$3217/B1 U$$1903/A2 U$$892/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1850/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _462_/CLK _325_/D VGND VGND VPWR VPWR _325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_256_ _267_/CLK _256_/D VGND VGND VPWR VPWR _256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_187_ _333_/CLK _187_/D VGND VGND VPWR VPWR _187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_63_5 dadda_fa_2_63_5/A dadda_fa_2_63_5/B dadda_fa_2_63_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_2/A dadda_fa_4_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater705 U$$56/A1 VGND VGND VPWR VPWR U$$4303/A1 sky130_fd_sc_hd__buf_12
Xrepeater716 _572_/Q VGND VGND VPWR VPWR U$$4156/B1 sky130_fd_sc_hd__buf_12
Xrepeater727 _567_/Q VGND VGND VPWR VPWR U$$38/A1 sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_1_clk _431_/CLK VGND VGND VPWR VPWR _429_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_56_4 dadda_fa_2_56_4/A dadda_fa_2_56_4/B dadda_fa_2_56_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/CIN dadda_fa_3_56_3/CIN sky130_fd_sc_hd__fa_1
XU$$4420 _566_/Q U$$4388/X _567_/Q U$$4389/X VGND VGND VPWR VPWR U$$4421/A sky130_fd_sc_hd__a22o_1
Xrepeater738 _562_/Q VGND VGND VPWR VPWR U$$28/A1 sky130_fd_sc_hd__buf_12
XFILLER_42_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater749 U$$4265/A1 VGND VGND VPWR VPWR U$$975/B1 sky130_fd_sc_hd__buf_12
XU$$4431 U$$4431/A U$$4431/B VGND VGND VPWR VPWR U$$4431/X sky130_fd_sc_hd__xor2_2
XU$$4442 U$$4442/A1 U$$4388/X _578_/Q U$$4389/X VGND VGND VPWR VPWR U$$4443/A sky130_fd_sc_hd__a22o_2
XU$$4453 U$$4453/A U$$4453/B VGND VGND VPWR VPWR U$$4453/X sky130_fd_sc_hd__xor2_4
XFILLER_93_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4464 U$$765/A1 U$$4388/X U$$82/A1 U$$4389/X VGND VGND VPWR VPWR U$$4465/A sky130_fd_sc_hd__a22o_2
XFILLER_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_49_3 dadda_fa_2_49_3/A dadda_fa_2_49_3/B dadda_fa_2_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/B dadda_fa_3_49_3/B sky130_fd_sc_hd__fa_1
XU$$4475 U$$4475/A U$$4475/B VGND VGND VPWR VPWR U$$4475/X sky130_fd_sc_hd__xor2_1
XU$$3730 U$$3730/A U$$3756/B VGND VGND VPWR VPWR U$$3730/X sky130_fd_sc_hd__xor2_1
XFILLER_53_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3741 U$$4289/A1 U$$3795/A2 U$$4289/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3742/A
+ sky130_fd_sc_hd__a22o_1
XU$$4486 U$$4486/A1 U$$4388/X U$$787/B1 U$$4389/X VGND VGND VPWR VPWR U$$4487/A sky130_fd_sc_hd__a22o_1
XU$$3752 U$$3752/A U$$3794/B VGND VGND VPWR VPWR U$$3752/X sky130_fd_sc_hd__xor2_1
XU$$4497 U$$4497/A U$$4497/B VGND VGND VPWR VPWR U$$4497/X sky130_fd_sc_hd__xor2_2
XFILLER_18_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3763 _580_/Q U$$3795/A2 _581_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3764/A sky130_fd_sc_hd__a22o_1
XU$$3774 U$$3774/A _671_/Q VGND VGND VPWR VPWR U$$3774/X sky130_fd_sc_hd__xor2_1
XU$$3785 U$$771/A1 U$$3703/X U$$771/B1 U$$3704/X VGND VGND VPWR VPWR U$$3786/A sky130_fd_sc_hd__a22o_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_19_1 dadda_fa_5_19_1/A dadda_fa_5_19_1/B dadda_fa_5_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/B dadda_fa_7_19_0/A sky130_fd_sc_hd__fa_1
XU$$3796 U$$3796/A _671_/Q VGND VGND VPWR VPWR U$$3796/X sky130_fd_sc_hd__xor2_1
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_3 U$$1306/X U$$1439/X U$$1572/X VGND VGND VPWR VPWR dadda_fa_2_52_1/B
+ dadda_fa_2_51_4/B sky130_fd_sc_hd__fa_1
XFILLER_83_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$907 U$$907/A U$$943/B VGND VGND VPWR VPWR U$$907/X sky130_fd_sc_hd__xor2_1
XU$$918 U$$96/A1 U$$928/A2 U$$96/B1 U$$928/B2 VGND VGND VPWR VPWR U$$919/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_2 U$$893/X U$$1026/X U$$1159/X VGND VGND VPWR VPWR dadda_fa_2_45_3/A
+ dadda_fa_2_44_5/A sky130_fd_sc_hd__fa_1
XU$$929 U$$929/A U$$943/B VGND VGND VPWR VPWR U$$929/X sky130_fd_sc_hd__xor2_1
XFILLER_56_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_21_1 dadda_fa_4_21_1/A dadda_fa_4_21_1/B dadda_fa_4_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/B dadda_fa_5_21_1/B sky130_fd_sc_hd__fa_2
XFILLER_55_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_14_0 U$$301/X U$$434/X U$$567/X VGND VGND VPWR VPWR dadda_fa_5_15_0/A
+ dadda_fa_5_14_1/A sky130_fd_sc_hd__fa_2
XFILLER_52_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_66_3 dadda_fa_3_66_3/A dadda_fa_3_66_3/B dadda_fa_3_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/B dadda_fa_4_66_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_59_2 dadda_fa_3_59_2/A dadda_fa_3_59_2/B dadda_fa_3_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/A dadda_fa_4_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3004 U$$3004/A U$$3004/B VGND VGND VPWR VPWR U$$3004/X sky130_fd_sc_hd__xor2_1
XU$$3015 _660_/Q VGND VGND VPWR VPWR U$$3017/B sky130_fd_sc_hd__inv_1
XFILLER_46_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_29_0 dadda_fa_6_29_0/A dadda_fa_6_29_0/B dadda_fa_6_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_30_0/B dadda_fa_7_29_0/CIN sky130_fd_sc_hd__fa_2
XU$$3026 U$$4122/A1 U$$3090/A2 U$$14/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3027/A sky130_fd_sc_hd__a22o_1
XU$$3037 U$$3037/A U$$3085/B VGND VGND VPWR VPWR U$$3037/X sky130_fd_sc_hd__xor2_1
XU$$3048 _565_/Q U$$3090/A2 U$$4283/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3049/A sky130_fd_sc_hd__a22o_1
XU$$2303 U$$2303/A U$$2327/B VGND VGND VPWR VPWR U$$2303/X sky130_fd_sc_hd__xor2_1
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3059 U$$3059/A U$$3085/B VGND VGND VPWR VPWR U$$3059/X sky130_fd_sc_hd__xor2_1
XU$$2314 _609_/Q U$$2326/A2 _610_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2315/A sky130_fd_sc_hd__a22o_1
XFILLER_189_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2325 U$$2325/A _649_/Q VGND VGND VPWR VPWR U$$2325/X sky130_fd_sc_hd__xor2_1
XFILLER_74_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2336 U$$2336/A U$$2432/B VGND VGND VPWR VPWR U$$2336/X sky130_fd_sc_hd__xor2_1
XU$$1602 U$$1602/A _639_/Q VGND VGND VPWR VPWR U$$1602/X sky130_fd_sc_hd__xor2_1
XU$$2347 U$$18/A1 U$$2333/X U$$20/A1 U$$2334/X VGND VGND VPWR VPWR U$$2348/A sky130_fd_sc_hd__a22o_1
XFILLER_188_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2358 U$$2358/A U$$2436/B VGND VGND VPWR VPWR U$$2358/X sky130_fd_sc_hd__xor2_1
XU$$1613 U$$654/A1 U$$1641/A2 U$$930/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1614/A sky130_fd_sc_hd__a22o_1
XU$$2369 U$$3191/A1 U$$2421/A2 U$$4289/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2370/A
+ sky130_fd_sc_hd__a22o_1
XU$$1624 U$$1624/A U$$1643/A VGND VGND VPWR VPWR U$$1624/X sky130_fd_sc_hd__xor2_1
XU$$1635 U$$950/A1 U$$1641/A2 U$$952/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1636/A sky130_fd_sc_hd__a22o_1
XU$$1646 U$$1781/A VGND VGND VPWR VPWR U$$1646/Y sky130_fd_sc_hd__inv_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1657 U$$1657/A U$$1727/B VGND VGND VPWR VPWR U$$1657/X sky130_fd_sc_hd__xor2_1
XU$$1668 U$$4271/A1 U$$1726/A2 U$$4273/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1669/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1679 U$$1679/A U$$1727/B VGND VGND VPWR VPWR U$$1679/X sky130_fd_sc_hd__xor2_1
XFILLER_148_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_308_ _463_/CLK _308_/D VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_239_ _500_/CLK _239_/D VGND VGND VPWR VPWR _239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_61_2 dadda_fa_2_61_2/A dadda_fa_2_61_2/B dadda_fa_2_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/A dadda_fa_3_61_3/A sky130_fd_sc_hd__fa_2
XFILLER_112_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater502 U$$1786/X VGND VGND VPWR VPWR U$$1867/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$309 final_adder.U$$308/A final_adder.U$$233/X final_adder.U$$235/X
+ VGND VGND VPWR VPWR final_adder.U$$309/X sky130_fd_sc_hd__a21o_1
Xrepeater513 U$$1101/X VGND VGND VPWR VPWR U$$1200/B2 sky130_fd_sc_hd__buf_12
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater524 _673_/Q VGND VGND VPWR VPWR U$$3969/B sky130_fd_sc_hd__buf_12
XFILLER_66_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_54_1 dadda_fa_2_54_1/A dadda_fa_2_54_1/B dadda_fa_2_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/CIN dadda_fa_3_54_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_78_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater535 _667_/Q VGND VGND VPWR VPWR U$$3536/B sky130_fd_sc_hd__buf_12
Xrepeater546 U$$2996/B VGND VGND VPWR VPWR U$$2960/B sky130_fd_sc_hd__buf_12
Xrepeater557 _653_/Q VGND VGND VPWR VPWR U$$2603/A sky130_fd_sc_hd__buf_12
XFILLER_133_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_31_0 dadda_fa_5_31_0/A dadda_fa_5_31_0/B dadda_fa_5_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/A dadda_fa_6_31_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater568 U$$2055/A VGND VGND VPWR VPWR U$$2023/B sky130_fd_sc_hd__buf_12
Xrepeater579 _639_/Q VGND VGND VPWR VPWR U$$1614/B sky130_fd_sc_hd__buf_12
XU$$4250 U$$4332/B U$$4250/B VGND VGND VPWR VPWR U$$4250/X sky130_fd_sc_hd__and2_1
Xdadda_fa_2_47_0 U$$2761/X U$$2894/X U$$3027/X VGND VGND VPWR VPWR dadda_fa_3_48_0/B
+ dadda_fa_3_47_2/B sky130_fd_sc_hd__fa_1
XU$$4261 _555_/Q U$$4381/A2 _556_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4262/A sky130_fd_sc_hd__a22o_1
XU$$4272 U$$4272/A _679_/Q VGND VGND VPWR VPWR U$$4272/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4283 U$$4283/A1 U$$4251/X U$$4285/A1 U$$4252/X VGND VGND VPWR VPWR U$$4284/A sky130_fd_sc_hd__a22o_1
XFILLER_168_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4294 U$$4294/A U$$4384/A VGND VGND VPWR VPWR U$$4294/X sky130_fd_sc_hd__xor2_2
XFILLER_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3560 U$$3560/A U$$3561/A VGND VGND VPWR VPWR U$$3560/X sky130_fd_sc_hd__xor2_1
XFILLER_37_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3571 U$$3571/A U$$3625/B VGND VGND VPWR VPWR U$$3571/X sky130_fd_sc_hd__xor2_1
XU$$3582 U$$979/A1 U$$3624/A2 U$$22/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3583/A sky130_fd_sc_hd__a22o_1
XU$$3593 U$$3593/A U$$3698/A VGND VGND VPWR VPWR U$$3593/X sky130_fd_sc_hd__xor2_1
XU$$2870 _613_/Q U$$2870/A2 _614_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2871/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_8_1 U$$623/B input245/X dadda_ha_4_8_0/SUM VGND VGND VPWR VPWR dadda_fa_6_9_0/B
+ dadda_fa_7_8_0/A sky130_fd_sc_hd__fa_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2881 U$$2879/Y _658_/Q _657_/Q U$$2880/X U$$2877/Y VGND VGND VPWR VPWR U$$2881/X
+ sky130_fd_sc_hd__a32o_4
XU$$2892 U$$2892/A U$$2996/B VGND VGND VPWR VPWR U$$2892/X sky130_fd_sc_hd__xor2_1
XFILLER_178_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_76_2 dadda_fa_4_76_2/A dadda_fa_4_76_2/B dadda_fa_4_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/CIN dadda_fa_5_76_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_69_1 dadda_fa_4_69_1/A dadda_fa_4_69_1/B dadda_fa_4_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/B dadda_fa_5_69_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_46_0 dadda_fa_7_46_0/A dadda_fa_7_46_0/B dadda_fa_7_46_0/CIN VGND VGND
+ VPWR VPWR _471_/D _342_/D sky130_fd_sc_hd__fa_1
XFILLER_130_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$704 U$$704/A U$$784/B VGND VGND VPWR VPWR U$$704/X sky130_fd_sc_hd__xor2_2
XFILLER_112_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$715 U$$28/B1 U$$817/A2 U$$32/A1 U$$785/B2 VGND VGND VPWR VPWR U$$716/A sky130_fd_sc_hd__a22o_1
X_590_ _601_/CLK _590_/D VGND VGND VPWR VPWR _590_/Q sky130_fd_sc_hd__dfxtp_4
XU$$726 U$$726/A U$$784/B VGND VGND VPWR VPWR U$$726/X sky130_fd_sc_hd__xor2_1
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$737 U$$50/B1 U$$785/A2 U$$876/A1 U$$785/B2 VGND VGND VPWR VPWR U$$738/A sky130_fd_sc_hd__a22o_1
XU$$748 U$$748/A U$$784/B VGND VGND VPWR VPWR U$$748/X sky130_fd_sc_hd__xor2_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$759 U$$759/A1 U$$817/A2 U$$759/B1 U$$817/B2 VGND VGND VPWR VPWR U$$760/A sky130_fd_sc_hd__a22o_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_71_1 dadda_fa_3_71_1/A dadda_fa_3_71_1/B dadda_fa_3_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/CIN dadda_fa_4_71_2/A sky130_fd_sc_hd__fa_2
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_64_0 dadda_fa_3_64_0/A dadda_fa_3_64_0/B dadda_fa_3_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/B dadda_fa_4_64_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2100 U$$2100/A U$$2118/B VGND VGND VPWR VPWR U$$2100/X sky130_fd_sc_hd__xor2_1
XU$$2111 U$$878/A1 U$$2117/A2 U$$4442/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2112/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_100_1 dadda_fa_4_100_1/A dadda_fa_4_100_1/B dadda_fa_4_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/B dadda_fa_5_100_1/B sky130_fd_sc_hd__fa_1
XU$$2122 U$$2122/A _647_/Q VGND VGND VPWR VPWR U$$2122/X sky130_fd_sc_hd__xor2_2
XU$$2133 U$$78/A1 U$$2059/X U$$765/A1 U$$2060/X VGND VGND VPWR VPWR U$$2134/A sky130_fd_sc_hd__a22o_1
XU$$2144 U$$2144/A _647_/Q VGND VGND VPWR VPWR U$$2144/X sky130_fd_sc_hd__xor2_1
XFILLER_23_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1410 U$$3191/A1 U$$1472/A2 U$$3876/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1411/A
+ sky130_fd_sc_hd__a22o_1
XU$$2155 _598_/Q U$$2161/A2 _599_/Q U$$2161/B2 VGND VGND VPWR VPWR U$$2156/A sky130_fd_sc_hd__a22o_1
XU$$1421 U$$1421/A U$$1479/B VGND VGND VPWR VPWR U$$1421/X sky130_fd_sc_hd__xor2_1
XU$$2166 U$$2166/A U$$2192/A VGND VGND VPWR VPWR U$$2166/X sky130_fd_sc_hd__xor2_1
XU$$2177 U$$944/A1 U$$2189/A2 U$$946/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2178/A sky130_fd_sc_hd__a22o_1
XU$$1432 U$$62/A1 U$$1472/A2 U$$64/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1433/A sky130_fd_sc_hd__a22o_1
XU$$1443 U$$1443/A U$$1505/B VGND VGND VPWR VPWR U$$1443/X sky130_fd_sc_hd__xor2_1
XU$$2188 U$$2188/A U$$2192/A VGND VGND VPWR VPWR U$$2188/X sky130_fd_sc_hd__xor2_1
XU$$2199 U$$2199/A U$$2289/B VGND VGND VPWR VPWR U$$2199/X sky130_fd_sc_hd__xor2_1
XU$$1454 U$$84/A1 U$$1472/A2 U$$908/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1455/A sky130_fd_sc_hd__a22o_1
XU$$1465 U$$1465/A U$$1479/B VGND VGND VPWR VPWR U$$1465/X sky130_fd_sc_hd__xor2_1
XFILLER_43_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1476 _601_/Q U$$1374/X U$$928/B1 U$$1375/X VGND VGND VPWR VPWR U$$1477/A sky130_fd_sc_hd__a22o_1
XFILLER_31_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_121_0 dadda_fa_7_121_0/A dadda_fa_7_121_0/B dadda_fa_7_121_0/CIN VGND
+ VGND VPWR VPWR _546_/D _417_/D sky130_fd_sc_hd__fa_2
XU$$1487 U$$1487/A U$$1505/B VGND VGND VPWR VPWR U$$1487/X sky130_fd_sc_hd__xor2_1
XFILLER_176_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1498 _612_/Q U$$1374/X U$$4514/A1 U$$1375/X VGND VGND VPWR VPWR U$$1499/A sky130_fd_sc_hd__a22o_1
XFILLER_188_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_86_1 dadda_fa_5_86_1/A dadda_fa_5_86_1/B dadda_fa_5_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/B dadda_fa_7_86_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_79_0 dadda_fa_5_79_0/A dadda_fa_5_79_0/B dadda_fa_5_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/A dadda_fa_6_79_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_144_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_78_8 U$$4419/X input232/X dadda_fa_1_78_8/CIN VGND VGND VPWR VPWR dadda_fa_2_79_3/A
+ dadda_fa_3_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_98_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$106 _530_/Q _402_/Q VGND VGND VPWR VPWR final_adder.U$$601/B1 final_adder.U$$728/A
+ sky130_fd_sc_hd__ha_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$117 _541_/Q _413_/Q VGND VGND VPWR VPWR final_adder.U$$245/B1 final_adder.U$$739/A
+ sky130_fd_sc_hd__ha_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$139 final_adder.U$$633/A final_adder.U$$505/B1 final_adder.U$$139/B1
+ VGND VGND VPWR VPWR final_adder.U$$139/X sky130_fd_sc_hd__a21o_1
XFILLER_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater387 U$$928/A2 VGND VGND VPWR VPWR U$$910/A2 sky130_fd_sc_hd__buf_12
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater398 U$$4114/X VGND VGND VPWR VPWR U$$4198/A2 sky130_fd_sc_hd__buf_12
XU$$4080 U$$4080/A U$$4109/A VGND VGND VPWR VPWR U$$4080/X sky130_fd_sc_hd__xor2_1
XFILLER_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4091 U$$4502/A1 U$$4107/A2 U$$4504/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3390 _599_/Q U$$3292/X _600_/Q U$$3293/X VGND VGND VPWR VPWR U$$3391/A sky130_fd_sc_hd__a22o_1
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_81_0 dadda_fa_4_81_0/A dadda_fa_4_81_0/B dadda_fa_4_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/A dadda_fa_5_81_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_102_3 dadda_fa_3_102_3/A dadda_fa_3_102_3/B dadda_fa_3_102_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/B dadda_fa_4_102_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput102 b[43] VGND VGND VPWR VPWR _595_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput113 b[53] VGND VGND VPWR VPWR _605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput124 b[63] VGND VGND VPWR VPWR _615_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput135 c[105] VGND VGND VPWR VPWR input135/X sky130_fd_sc_hd__buf_2
Xinput146 c[115] VGND VGND VPWR VPWR input146/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput157 c[125] VGND VGND VPWR VPWR input157/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput168 c[1] VGND VGND VPWR VPWR input168/X sky130_fd_sc_hd__buf_4
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$640 final_adder.U$$640/A final_adder.U$$640/B VGND VGND VPWR VPWR
+ _186_/D sky130_fd_sc_hd__xor2_2
Xinput179 c[2] VGND VGND VPWR VPWR input179/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$651 final_adder.U$$651/A final_adder.U$$651/B VGND VGND VPWR VPWR
+ _197_/D sky130_fd_sc_hd__xor2_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_642_ _642_/CLK _642_/D VGND VGND VPWR VPWR _642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$662 final_adder.U$$662/A final_adder.U$$662/B VGND VGND VPWR VPWR
+ _208_/D sky130_fd_sc_hd__xor2_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$501 U$$90/A1 U$$545/A2 U$$92/A1 U$$416/X VGND VGND VPWR VPWR U$$502/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_109_0 dadda_fa_6_109_0/A dadda_fa_6_109_0/B dadda_fa_6_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_110_0/B dadda_fa_7_109_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$673 final_adder.U$$673/A final_adder.U$$673/B VGND VGND VPWR VPWR
+ _219_/D sky130_fd_sc_hd__xor2_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$512 U$$512/A U$$547/A VGND VGND VPWR VPWR U$$512/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$684 final_adder.U$$684/A final_adder.U$$684/B VGND VGND VPWR VPWR
+ _230_/D sky130_fd_sc_hd__xor2_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$523 U$$934/A1 U$$545/A2 U$$799/A1 U$$416/X VGND VGND VPWR VPWR U$$524/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$695 final_adder.U$$695/A final_adder.U$$695/B VGND VGND VPWR VPWR
+ _241_/D sky130_fd_sc_hd__xor2_1
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$534 U$$534/A _623_/Q VGND VGND VPWR VPWR U$$534/X sky130_fd_sc_hd__xor2_1
XFILLER_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$545 U$$956/A1 U$$545/A2 U$$545/B1 U$$416/X VGND VGND VPWR VPWR U$$546/A sky130_fd_sc_hd__a22o_1
XFILLER_72_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_573_ _573_/CLK _573_/D VGND VGND VPWR VPWR _573_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$556 _552_/Q U$$626/A2 U$$969/A1 U$$553/X VGND VGND VPWR VPWR U$$557/A sky130_fd_sc_hd__a22o_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_3 dadda_fa_3_29_3/A dadda_fa_3_29_3/B dadda_fa_3_29_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/B dadda_fa_4_29_2/CIN sky130_fd_sc_hd__fa_1
XU$$567 U$$567/A U$$623/B VGND VGND VPWR VPWR U$$567/X sky130_fd_sc_hd__xor2_1
XFILLER_60_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$578 U$$28/B1 U$$626/A2 U$$32/A1 U$$553/X VGND VGND VPWR VPWR U$$579/A sky130_fd_sc_hd__a22o_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$589 U$$589/A U$$623/B VGND VGND VPWR VPWR U$$589/X sky130_fd_sc_hd__xor2_1
XFILLER_25_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_96_0 dadda_fa_6_96_0/A dadda_fa_6_96_0/B dadda_fa_6_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_97_0/B dadda_fa_7_96_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_184_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_2_32_5 U$$2066/X U$$2199/X VGND VGND VPWR VPWR dadda_fa_3_33_2/A dadda_fa_4_32_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_31_3 U$$1266/X U$$1399/X U$$1532/X VGND VGND VPWR VPWR dadda_fa_3_32_1/CIN
+ dadda_fa_3_31_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1240 U$$1240/A U$$1336/B VGND VGND VPWR VPWR U$$1240/X sky130_fd_sc_hd__xor2_1
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1251 U$$18/A1 U$$1237/X U$$20/A1 U$$1238/X VGND VGND VPWR VPWR U$$1252/A sky130_fd_sc_hd__a22o_1
XU$$1262 U$$1262/A U$$1336/B VGND VGND VPWR VPWR U$$1262/X sky130_fd_sc_hd__xor2_1
XU$$1273 U$$3191/A1 U$$1341/A2 U$$3876/B1 U$$1341/B2 VGND VGND VPWR VPWR U$$1274/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1284 U$$1284/A U$$1342/B VGND VGND VPWR VPWR U$$1284/X sky130_fd_sc_hd__xor2_1
XU$$1295 U$$62/A1 U$$1341/A2 U$$64/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1296/A sky130_fd_sc_hd__a22o_1
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_6 U$$3764/X U$$3897/X U$$4030/X VGND VGND VPWR VPWR dadda_fa_2_84_3/CIN
+ dadda_fa_3_83_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_76_5 U$$3484/X U$$3617/X U$$3750/X VGND VGND VPWR VPWR dadda_fa_2_77_2/A
+ dadda_fa_2_76_5/A sky130_fd_sc_hd__fa_1
XFILLER_98_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_4 U$$4002/X U$$4135/X U$$4268/X VGND VGND VPWR VPWR dadda_fa_2_70_1/CIN
+ dadda_fa_2_69_4/CIN sky130_fd_sc_hd__fa_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_39_2 dadda_fa_4_39_2/A dadda_fa_4_39_2/B dadda_fa_4_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/CIN dadda_fa_5_39_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_100_0 U$$4330/X U$$4463/X input130/X VGND VGND VPWR VPWR dadda_fa_4_101_0/B
+ dadda_fa_4_100_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_123_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_64_3 U$$1332/X U$$1465/X U$$1598/X VGND VGND VPWR VPWR dadda_fa_1_65_6/B
+ dadda_fa_1_64_8/B sky130_fd_sc_hd__fa_2
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_41_2 dadda_fa_3_41_2/A dadda_fa_3_41_2/B dadda_fa_3_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/A dadda_fa_4_41_2/B sky130_fd_sc_hd__fa_2
XFILLER_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$481 final_adder.U$$304/B final_adder.U$$718/B final_adder.U$$225/X
+ VGND VGND VPWR VPWR final_adder.U$$720/B sky130_fd_sc_hd__a21o_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_625_ _642_/CLK _625_/D VGND VGND VPWR VPWR _625_/Q sky130_fd_sc_hd__dfxtp_4
XU$$320 U$$46/A1 U$$278/X _572_/Q U$$279/X VGND VGND VPWR VPWR U$$321/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_1 dadda_fa_3_34_1/A dadda_fa_3_34_1/B dadda_fa_3_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/CIN dadda_fa_4_34_2/A sky130_fd_sc_hd__fa_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$331 U$$331/A U$$391/B VGND VGND VPWR VPWR U$$331/X sky130_fd_sc_hd__xor2_1
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$342 U$$68/A1 U$$278/X U$$68/B1 U$$279/X VGND VGND VPWR VPWR U$$343/A sky130_fd_sc_hd__a22o_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$353 U$$353/A U$$391/B VGND VGND VPWR VPWR U$$353/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_11_0 dadda_fa_6_11_0/A dadda_fa_6_11_0/B dadda_fa_6_11_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_12_0/B dadda_fa_7_11_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_72_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_27_0 U$$1125/X U$$1258/X U$$1391/X VGND VGND VPWR VPWR dadda_fa_4_28_0/B
+ dadda_fa_4_27_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$364 U$$90/A1 U$$278/X U$$92/A1 U$$279/X VGND VGND VPWR VPWR U$$365/A sky130_fd_sc_hd__a22o_1
XU$$375 U$$375/A U$$391/B VGND VGND VPWR VPWR U$$375/X sky130_fd_sc_hd__xor2_1
X_556_ _649_/CLK _556_/D VGND VGND VPWR VPWR _556_/Q sky130_fd_sc_hd__dfxtp_4
XU$$386 U$$934/A1 U$$278/X U$$799/A1 U$$279/X VGND VGND VPWR VPWR U$$387/A sky130_fd_sc_hd__a22o_1
XU$$397 U$$397/A _621_/Q VGND VGND VPWR VPWR U$$397/X sky130_fd_sc_hd__xor2_1
X_487_ _490_/CLK _487_/D VGND VGND VPWR VPWR _487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_93_5 dadda_fa_2_93_5/A dadda_fa_2_93_5/B dadda_fa_2_93_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_94_2/A dadda_fa_4_93_0/A sky130_fd_sc_hd__fa_2
XFILLER_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_86_4 dadda_fa_2_86_4/A dadda_fa_2_86_4/B dadda_fa_2_86_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/CIN dadda_fa_3_86_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_126_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_79_3 dadda_fa_2_79_3/A dadda_fa_2_79_3/B dadda_fa_2_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/B dadda_fa_3_79_3/B sky130_fd_sc_hd__fa_2
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_49_1 dadda_fa_5_49_1/A dadda_fa_5_49_1/B dadda_fa_5_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/B dadda_fa_7_49_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_746__798 VGND VGND VPWR VPWR _746__798/HI U$$3157/A1 sky130_fd_sc_hd__conb_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_102_2 U$$3403/X U$$3536/X U$$3669/X VGND VGND VPWR VPWR dadda_fa_3_103_2/CIN
+ dadda_fa_3_102_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1070 U$$1070/A U$$998/B VGND VGND VPWR VPWR U$$1070/X sky130_fd_sc_hd__xor2_1
XFILLER_189_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1081 U$$944/A1 U$$963/X U$$946/A1 U$$964/X VGND VGND VPWR VPWR U$$1082/A sky130_fd_sc_hd__a22o_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1092 U$$1092/A _631_/Q VGND VGND VPWR VPWR U$$1092/X sky130_fd_sc_hd__xor2_1
XFILLER_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_123_1 U$$4509/X input155/X dadda_fa_5_123_1/CIN VGND VGND VPWR VPWR dadda_fa_6_124_0/B
+ dadda_fa_7_123_0/A sky130_fd_sc_hd__fa_1
XFILLER_13_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_116_0 dadda_fa_5_116_0/A dadda_fa_5_116_0/B dadda_fa_5_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/A dadda_fa_6_116_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_81_3 U$$2430/X U$$2563/X U$$2696/X VGND VGND VPWR VPWR dadda_fa_2_82_2/A
+ dadda_fa_2_81_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_74_2 U$$2549/X U$$2682/X U$$2815/X VGND VGND VPWR VPWR dadda_fa_2_75_1/A
+ dadda_fa_2_74_4/A sky130_fd_sc_hd__fa_1
XFILLER_99_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_51_1 dadda_fa_4_51_1/A dadda_fa_4_51_1/B dadda_fa_4_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/B dadda_fa_5_51_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_1 U$$2934/X U$$3067/X U$$3200/X VGND VGND VPWR VPWR dadda_fa_2_68_0/CIN
+ dadda_fa_2_67_3/CIN sky130_fd_sc_hd__fa_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_44_0 dadda_fa_4_44_0/A dadda_fa_4_44_0/B dadda_fa_4_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/A dadda_fa_5_44_1/A sky130_fd_sc_hd__fa_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _543_/CLK _410_/D VGND VGND VPWR VPWR _410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ _469_/CLK _341_/D VGND VGND VPWR VPWR _341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_695__915 VGND VGND VPWR VPWR _695__915/HI _695__915/LO sky130_fd_sc_hd__conb_1
XFILLER_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ _280_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_96_3 dadda_fa_3_96_3/A dadda_fa_3_96_3/B dadda_fa_3_96_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/B dadda_fa_4_96_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_89_2 dadda_fa_3_89_2/A dadda_fa_3_89_2/B dadda_fa_3_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/A dadda_fa_4_89_2/B sky130_fd_sc_hd__fa_2
XFILLER_108_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_59_0 dadda_fa_6_59_0/A dadda_fa_6_59_0/B dadda_fa_6_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_60_0/B dadda_fa_7_59_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_62_0 U$$131/X U$$264/X U$$397/X VGND VGND VPWR VPWR dadda_fa_1_63_5/B
+ dadda_fa_1_62_7/B sky130_fd_sc_hd__fa_1
XFILLER_65_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3901 U$$3901/A U$$3929/B VGND VGND VPWR VPWR U$$3901/X sky130_fd_sc_hd__xor2_1
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3912 U$$76/A1 U$$3912/A2 _587_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3913/A sky130_fd_sc_hd__a22o_1
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3923 U$$3923/A _673_/Q VGND VGND VPWR VPWR U$$3923/X sky130_fd_sc_hd__xor2_1
XFILLER_18_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3934 U$$98/A1 U$$3970/A2 U$$98/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3935/A sky130_fd_sc_hd__a22o_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3945 U$$3945/A _673_/Q VGND VGND VPWR VPWR U$$3945/X sky130_fd_sc_hd__xor2_1
XU$$3956 U$$4504/A1 U$$3970/A2 U$$4506/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3957/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3967 U$$3967/A U$$3969/B VGND VGND VPWR VPWR U$$3967/X sky130_fd_sc_hd__xor2_1
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3978 U$$3976/B _673_/Q _674_/Q U$$3973/Y VGND VGND VPWR VPWR U$$3978/X sky130_fd_sc_hd__a22o_4
X_608_ _611_/CLK _608_/D VGND VGND VPWR VPWR _608_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$150 U$$150/A U$$242/B VGND VGND VPWR VPWR U$$150/X sky130_fd_sc_hd__xor2_1
XU$$3989 _556_/Q U$$3977/X U$$975/B1 U$$3978/X VGND VGND VPWR VPWR U$$3990/A sky130_fd_sc_hd__a22o_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$161 _560_/Q U$$141/X U$$26/A1 U$$142/X VGND VGND VPWR VPWR U$$162/A sky130_fd_sc_hd__a22o_1
XFILLER_73_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$172 U$$172/A U$$262/B VGND VGND VPWR VPWR U$$172/X sky130_fd_sc_hd__xor2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$183 U$$46/A1 U$$141/X U$$48/A1 U$$142/X VGND VGND VPWR VPWR U$$184/A sky130_fd_sc_hd__a22o_1
XU$$194 U$$194/A U$$262/B VGND VGND VPWR VPWR U$$194/X sky130_fd_sc_hd__xor2_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_539_ _543_/CLK _539_/D VGND VGND VPWR VPWR _539_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_91_2 U$$3913/X U$$4046/X U$$4179/X VGND VGND VPWR VPWR dadda_fa_3_92_1/A
+ dadda_fa_3_91_3/A sky130_fd_sc_hd__fa_1
XFILLER_127_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_84_1 U$$4431/X input239/X dadda_fa_2_84_1/CIN VGND VGND VPWR VPWR dadda_fa_3_85_0/CIN
+ dadda_fa_3_84_2/CIN sky130_fd_sc_hd__fa_2
Xoutput258 _268_/Q VGND VGND VPWR VPWR o[100] sky130_fd_sc_hd__buf_2
Xoutput269 _278_/Q VGND VGND VPWR VPWR o[110] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_61_0 dadda_fa_5_61_0/A dadda_fa_5_61_0/B dadda_fa_5_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/A dadda_fa_6_61_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_77_0 dadda_fa_2_77_0/A dadda_fa_2_77_0/B dadda_fa_2_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/B dadda_fa_3_77_2/B sky130_fd_sc_hd__fa_2
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_60_8 dadda_fa_1_60_8/A dadda_fa_1_60_8/B dadda_fa_1_60_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_3/A dadda_fa_3_60_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_53_7 U$$3172/X U$$3305/X U$$3438/X VGND VGND VPWR VPWR dadda_fa_2_54_2/CIN
+ dadda_fa_2_53_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_99_1 dadda_fa_4_99_1/A dadda_fa_4_99_1/B dadda_fa_4_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/B dadda_fa_5_99_1/B sky130_fd_sc_hd__fa_1
XFILLER_191_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_76_0 dadda_fa_7_76_0/A dadda_fa_7_76_0/B dadda_fa_7_76_0/CIN VGND VGND
+ VPWR VPWR _501_/D _372_/D sky130_fd_sc_hd__fa_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3208 U$$3208/A U$$3244/B VGND VGND VPWR VPWR U$$3208/X sky130_fd_sc_hd__xor2_1
XFILLER_19_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3219 U$$4178/A1 U$$3243/A2 U$$892/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3220/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2507 U$$2507/A U$$2533/B VGND VGND VPWR VPWR U$$2507/X sky130_fd_sc_hd__xor2_1
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2518 U$$50/B1 U$$2584/A2 U$$4438/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2519/A sky130_fd_sc_hd__a22o_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2529 U$$2529/A U$$2533/B VGND VGND VPWR VPWR U$$2529/X sky130_fd_sc_hd__xor2_1
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1806 U$$1806/A U$$1856/B VGND VGND VPWR VPWR U$$1806/X sky130_fd_sc_hd__xor2_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1817 U$$36/A1 U$$1867/A2 U$$38/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1818/A sky130_fd_sc_hd__a22o_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1828 U$$1828/A U$$1872/B VGND VGND VPWR VPWR U$$1828/X sky130_fd_sc_hd__xor2_1
XU$$1839 U$$880/A1 U$$1903/A2 U$$4170/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1840/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _458_/CLK _324_/D VGND VGND VPWR VPWR _324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_255_ _503_/CLK _255_/D VGND VGND VPWR VPWR _255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_186_ _333_/CLK _186_/D VGND VGND VPWR VPWR _186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_94_0 dadda_fa_3_94_0/A dadda_fa_3_94_0/B dadda_fa_3_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/B dadda_fa_4_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater706 _576_/Q VGND VGND VPWR VPWR U$$56/A1 sky130_fd_sc_hd__buf_12
Xrepeater717 U$$46/A1 VGND VGND VPWR VPWR U$$868/A1 sky130_fd_sc_hd__buf_12
Xrepeater728 _567_/Q VGND VGND VPWR VPWR U$$4285/A1 sky130_fd_sc_hd__buf_12
XU$$4410 _561_/Q U$$4388/X _562_/Q U$$4389/X VGND VGND VPWR VPWR U$$4411/A sky130_fd_sc_hd__a22o_1
XU$$4421 U$$4421/A U$$4421/B VGND VGND VPWR VPWR U$$4421/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_56_5 dadda_fa_2_56_5/A dadda_fa_2_56_5/B dadda_fa_2_56_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_2/A dadda_fa_4_56_0/A sky130_fd_sc_hd__fa_2
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater739 _561_/Q VGND VGND VPWR VPWR U$$26/A1 sky130_fd_sc_hd__buf_12
XU$$4432 _572_/Q U$$4388/X U$$735/A1 U$$4389/X VGND VGND VPWR VPWR U$$4433/A sky130_fd_sc_hd__a22o_1
XU$$4443 U$$4443/A U$$4443/B VGND VGND VPWR VPWR U$$4443/X sky130_fd_sc_hd__xor2_4
XU$$4454 U$$70/A1 U$$4388/X U$$70/B1 U$$4389/X VGND VGND VPWR VPWR U$$4455/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_4 dadda_fa_2_49_4/A dadda_fa_2_49_4/B dadda_fa_2_49_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/CIN dadda_fa_3_49_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4465 U$$4465/A U$$4465/B VGND VGND VPWR VPWR U$$4465/X sky130_fd_sc_hd__xor2_4
XU$$3720 U$$3720/A U$$3756/B VGND VGND VPWR VPWR U$$3720/X sky130_fd_sc_hd__xor2_1
XU$$4476 U$$4476/A1 U$$4388/X U$$94/A1 U$$4389/X VGND VGND VPWR VPWR U$$4477/A sky130_fd_sc_hd__a22o_1
XU$$3731 _564_/Q U$$3783/A2 _565_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3732/A sky130_fd_sc_hd__a22o_1
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3742 U$$3742/A U$$3794/B VGND VGND VPWR VPWR U$$3742/X sky130_fd_sc_hd__xor2_1
XU$$4487 U$$4487/A U$$4487/B VGND VGND VPWR VPWR U$$4487/X sky130_fd_sc_hd__xor2_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3753 _575_/Q U$$3795/A2 U$$4303/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3754/A sky130_fd_sc_hd__a22o_1
XU$$4498 U$$936/A1 U$$4388/X U$$4500/A1 U$$4389/X VGND VGND VPWR VPWR U$$4499/A sky130_fd_sc_hd__a22o_1
XU$$3764 U$$3764/A U$$3794/B VGND VGND VPWR VPWR U$$3764/X sky130_fd_sc_hd__xor2_1
XU$$3775 _586_/Q U$$3795/A2 _587_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3776/A sky130_fd_sc_hd__a22o_1
XFILLER_18_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3786 U$$3786/A U$$3835/A VGND VGND VPWR VPWR U$$3786/X sky130_fd_sc_hd__xor2_1
XFILLER_46_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3797 U$$98/A1 U$$3703/X U$$4484/A1 U$$3704/X VGND VGND VPWR VPWR U$$3798/A sky130_fd_sc_hd__a22o_1
XFILLER_61_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_1_45_5 U$$2092/X U$$2225/X VGND VGND VPWR VPWR dadda_fa_2_46_3/CIN dadda_fa_3_45_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_51_4 U$$1705/X U$$1838/X U$$1971/X VGND VGND VPWR VPWR dadda_fa_2_52_1/CIN
+ dadda_fa_2_51_4/CIN sky130_fd_sc_hd__fa_1
X_761__813 VGND VGND VPWR VPWR _761__813/HI U$$4107/B1 sky130_fd_sc_hd__conb_1
XFILLER_141_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$908 U$$908/A1 U$$928/A2 U$$88/A1 U$$928/B2 VGND VGND VPWR VPWR U$$909/A sky130_fd_sc_hd__a22o_1
XFILLER_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$919 U$$919/A U$$943/B VGND VGND VPWR VPWR U$$919/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_3 U$$1292/X U$$1425/X U$$1558/X VGND VGND VPWR VPWR dadda_fa_2_45_3/B
+ dadda_fa_2_44_5/B sky130_fd_sc_hd__fa_2
XFILLER_84_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_21_2 dadda_fa_4_21_2/A dadda_fa_4_21_2/B dadda_ha_3_21_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/CIN dadda_fa_5_21_1/CIN sky130_fd_sc_hd__fa_1
X_802__854 VGND VGND VPWR VPWR _802__854/HI U$$4449/B sky130_fd_sc_hd__conb_1
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_14_1 U$$700/X U$$833/X U$$966/X VGND VGND VPWR VPWR dadda_fa_5_15_0/B
+ dadda_fa_5_14_1/B sky130_fd_sc_hd__fa_1
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_59_3 dadda_fa_3_59_3/A dadda_fa_3_59_3/B dadda_fa_3_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/B dadda_fa_4_59_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3005 U$$950/A1 U$$3009/A2 U$$4514/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$3006/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3016 _661_/Q VGND VGND VPWR VPWR U$$3016/Y sky130_fd_sc_hd__inv_1
XFILLER_19_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3027 U$$3027/A U$$3085/B VGND VGND VPWR VPWR U$$3027/X sky130_fd_sc_hd__xor2_1
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3038 U$$4271/A1 U$$3090/A2 U$$4273/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3039/A
+ sky130_fd_sc_hd__a22o_1
XU$$3049 U$$3049/A U$$3109/B VGND VGND VPWR VPWR U$$3049/X sky130_fd_sc_hd__xor2_1
XFILLER_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2304 U$$4496/A1 U$$2326/A2 _605_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2305/A sky130_fd_sc_hd__a22o_1
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2315 U$$2315/A U$$2327/B VGND VGND VPWR VPWR U$$2315/X sky130_fd_sc_hd__xor2_1
XU$$2326 _615_/Q U$$2326/A2 U$$2326/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2327/A sky130_fd_sc_hd__a22o_1
XFILLER_90_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2337 U$$8/A1 U$$2333/X U$$8/B1 U$$2334/X VGND VGND VPWR VPWR U$$2338/A sky130_fd_sc_hd__a22o_1
XU$$2348 U$$2348/A U$$2432/B VGND VGND VPWR VPWR U$$2348/X sky130_fd_sc_hd__xor2_1
XU$$1603 U$$96/A1 U$$1605/A2 U$$96/B1 U$$1605/B2 VGND VGND VPWR VPWR U$$1604/A sky130_fd_sc_hd__a22o_1
XFILLER_90_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1614 U$$1614/A U$$1614/B VGND VGND VPWR VPWR U$$1614/X sky130_fd_sc_hd__xor2_1
XFILLER_90_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2359 U$$30/A1 U$$2421/A2 U$$30/B1 U$$2421/B2 VGND VGND VPWR VPWR U$$2360/A sky130_fd_sc_hd__a22o_1
XU$$1625 _607_/Q U$$1641/A2 _608_/Q U$$1641/B2 VGND VGND VPWR VPWR U$$1626/A sky130_fd_sc_hd__a22o_1
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1636 U$$1636/A _639_/Q VGND VGND VPWR VPWR U$$1636/X sky130_fd_sc_hd__xor2_1
XU$$1647 U$$1781/A U$$1647/B VGND VGND VPWR VPWR U$$1647/X sky130_fd_sc_hd__and2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1658 U$$12/B1 U$$1734/A2 U$$16/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1659/A sky130_fd_sc_hd__a22o_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1669 U$$1669/A U$$1739/B VGND VGND VPWR VPWR U$$1669/X sky130_fd_sc_hd__xor2_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_307_ _465_/CLK _307_/D VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_238_ _499_/CLK _238_/D VGND VGND VPWR VPWR _238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ _448_/CLK _169_/D VGND VGND VPWR VPWR _169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_3 dadda_fa_2_61_3/A dadda_fa_2_61_3/B dadda_fa_2_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/B dadda_fa_3_61_3/B sky130_fd_sc_hd__fa_1
Xrepeater503 U$$1770/B2 VGND VGND VPWR VPWR U$$1726/B2 sky130_fd_sc_hd__buf_12
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater514 U$$1101/X VGND VGND VPWR VPWR U$$1218/B2 sky130_fd_sc_hd__buf_12
Xrepeater525 _673_/Q VGND VGND VPWR VPWR U$$3893/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_54_2 dadda_fa_2_54_2/A dadda_fa_2_54_2/B dadda_fa_2_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/A dadda_fa_3_54_3/A sky130_fd_sc_hd__fa_2
Xrepeater536 _665_/Q VGND VGND VPWR VPWR U$$3413/B sky130_fd_sc_hd__buf_12
XFILLER_111_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater547 _659_/Q VGND VGND VPWR VPWR U$$2996/B sky130_fd_sc_hd__buf_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_31_1 dadda_fa_5_31_1/A dadda_fa_5_31_1/B dadda_fa_5_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/B dadda_fa_7_31_0/A sky130_fd_sc_hd__fa_1
XU$$4240 _613_/Q U$$4244/A2 U$$4379/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4241/A sky130_fd_sc_hd__a22o_1
Xrepeater558 _651_/Q VGND VGND VPWR VPWR U$$2432/B sky130_fd_sc_hd__buf_12
Xrepeater569 U$$2055/A VGND VGND VPWR VPWR U$$2021/B sky130_fd_sc_hd__buf_12
XFILLER_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4251 U$$4249/Y _678_/Q U$$4247/A U$$4250/X U$$4247/Y VGND VGND VPWR VPWR U$$4251/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_133_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4262 U$$4262/A _679_/Q VGND VGND VPWR VPWR U$$4262/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_47_1 U$$3160/X input198/X dadda_fa_2_47_1/CIN VGND VGND VPWR VPWR dadda_fa_3_48_0/CIN
+ dadda_fa_3_47_2/CIN sky130_fd_sc_hd__fa_2
XU$$4273 U$$4273/A1 U$$4251/X _562_/Q U$$4252/X VGND VGND VPWR VPWR U$$4274/A sky130_fd_sc_hd__a22o_1
XU$$4284 U$$4284/A U$$4332/B VGND VGND VPWR VPWR U$$4284/X sky130_fd_sc_hd__xor2_1
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_24_0 dadda_fa_5_24_0/A dadda_fa_5_24_0/B dadda_fa_5_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/A dadda_fa_6_24_0/CIN sky130_fd_sc_hd__fa_2
XU$$3550 U$$3550/A U$$3561/A VGND VGND VPWR VPWR U$$3550/X sky130_fd_sc_hd__xor2_1
XU$$4295 _572_/Q U$$4381/A2 U$$735/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4296/A sky130_fd_sc_hd__a22o_1
XFILLER_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3561 U$$3561/A VGND VGND VPWR VPWR U$$3561/Y sky130_fd_sc_hd__inv_1
XU$$3572 _553_/Q U$$3624/A2 U$$4122/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3573/A sky130_fd_sc_hd__a22o_1
XFILLER_19_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3583 U$$3583/A U$$3625/B VGND VGND VPWR VPWR U$$3583/X sky130_fd_sc_hd__xor2_1
XU$$3594 _564_/Q U$$3678/A2 _565_/Q U$$3678/B2 VGND VGND VPWR VPWR U$$3595/A sky130_fd_sc_hd__a22o_1
XU$$2860 U$$942/A1 U$$2744/X U$$4506/A1 U$$2745/X VGND VGND VPWR VPWR U$$2861/A sky130_fd_sc_hd__a22o_1
XU$$2871 U$$2871/A U$$2871/B VGND VGND VPWR VPWR U$$2871/X sky130_fd_sc_hd__xor2_1
XFILLER_34_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2882 U$$2880/B _657_/Q _658_/Q U$$2877/Y VGND VGND VPWR VPWR U$$2882/X sky130_fd_sc_hd__a22o_4
XU$$2893 U$$14/B1 U$$3009/A2 U$$4265/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2894/A sky130_fd_sc_hd__a22o_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_69_2 dadda_fa_4_69_2/A dadda_fa_4_69_2/B dadda_fa_4_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/CIN dadda_fa_5_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_1_36_1 U$$478/X U$$611/X VGND VGND VPWR VPWR dadda_fa_2_37_5/B dadda_fa_3_36_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_112_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_39_0 dadda_fa_7_39_0/A dadda_fa_7_39_0/B dadda_fa_7_39_0/CIN VGND VGND
+ VPWR VPWR _464_/D _335_/D sky130_fd_sc_hd__fa_1
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$705 U$$842/A1 U$$689/X U$$22/A1 U$$817/B2 VGND VGND VPWR VPWR U$$706/A sky130_fd_sc_hd__a22o_1
XFILLER_72_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$716 U$$716/A U$$784/B VGND VGND VPWR VPWR U$$716/X sky130_fd_sc_hd__xor2_1
XU$$727 _569_/Q U$$689/X _570_/Q U$$817/B2 VGND VGND VPWR VPWR U$$728/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_0 U$$91/X U$$224/X U$$357/X VGND VGND VPWR VPWR dadda_fa_2_43_3/A dadda_fa_2_42_4/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$738 U$$738/A U$$778/B VGND VGND VPWR VPWR U$$738/X sky130_fd_sc_hd__xor2_1
XFILLER_56_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$749 U$$64/A1 U$$785/A2 U$$66/A1 U$$785/B2 VGND VGND VPWR VPWR U$$750/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_71_2 dadda_fa_3_71_2/A dadda_fa_3_71_2/B dadda_fa_3_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/A dadda_fa_4_71_2/B sky130_fd_sc_hd__fa_2
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_64_1 dadda_fa_3_64_1/A dadda_fa_3_64_1/B dadda_fa_3_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/CIN dadda_fa_4_64_2/A sky130_fd_sc_hd__fa_1
XFILLER_126_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_41_0 dadda_fa_6_41_0/A dadda_fa_6_41_0/B dadda_fa_6_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_42_0/B dadda_fa_7_41_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_57_0 dadda_fa_3_57_0/A dadda_fa_3_57_0/B dadda_fa_3_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/B dadda_fa_4_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2101 U$$4291/B1 U$$2117/A2 U$$4156/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2102/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2112 U$$2112/A U$$2118/B VGND VGND VPWR VPWR U$$2112/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_100_2 dadda_fa_4_100_2/A dadda_fa_4_100_2/B dadda_fa_4_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/CIN dadda_fa_5_100_1/CIN sky130_fd_sc_hd__fa_1
XU$$2123 U$$3217/B1 U$$2161/A2 U$$892/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2124/A
+ sky130_fd_sc_hd__a22o_1
XU$$2134 U$$2134/A U$$2186/B VGND VGND VPWR VPWR U$$2134/X sky130_fd_sc_hd__xor2_1
XU$$2145 _593_/Q U$$2161/A2 U$$914/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2146/A sky130_fd_sc_hd__a22o_1
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1400 U$$28/B1 U$$1474/A2 U$$30/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1401/A sky130_fd_sc_hd__a22o_1
XU$$2156 U$$2156/A _647_/Q VGND VGND VPWR VPWR U$$2156/X sky130_fd_sc_hd__xor2_1
XU$$1411 U$$1411/A U$$1461/B VGND VGND VPWR VPWR U$$1411/X sky130_fd_sc_hd__xor2_1
XU$$2167 _604_/Q U$$2189/A2 U$$799/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2168/A sky130_fd_sc_hd__a22o_1
XFILLER_62_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1422 U$$50/B1 U$$1472/A2 U$$876/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1423/A sky130_fd_sc_hd__a22o_1
XU$$1433 U$$1433/A U$$1461/B VGND VGND VPWR VPWR U$$1433/X sky130_fd_sc_hd__xor2_1
XU$$2178 U$$2178/A U$$2192/A VGND VGND VPWR VPWR U$$2178/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2189 U$$956/A1 U$$2189/A2 U$$2189/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2190/A
+ sky130_fd_sc_hd__a22o_1
XU$$1444 U$$74/A1 U$$1472/A2 U$$2953/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1445/A sky130_fd_sc_hd__a22o_1
XU$$1455 U$$1455/A U$$1505/B VGND VGND VPWR VPWR U$$1455/X sky130_fd_sc_hd__xor2_1
XU$$1466 U$$94/B1 U$$1474/A2 U$$98/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1467/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1477 U$$1477/A U$$1505/B VGND VGND VPWR VPWR U$$1477/X sky130_fd_sc_hd__xor2_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1488 U$$940/A1 U$$1374/X U$$942/A1 U$$1375/X VGND VGND VPWR VPWR U$$1489/A sky130_fd_sc_hd__a22o_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1499 U$$1499/A U$$1505/B VGND VGND VPWR VPWR U$$1499/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_114_0 dadda_fa_7_114_0/A dadda_fa_7_114_0/B dadda_fa_7_114_0/CIN VGND
+ VGND VPWR VPWR _539_/D _410_/D sky130_fd_sc_hd__fa_2
XFILLER_184_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_79_1 dadda_fa_5_79_1/A dadda_fa_5_79_1/B dadda_fa_5_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/B dadda_fa_7_79_0/A sky130_fd_sc_hd__fa_1
XFILLER_171_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$107 _531_/Q _403_/Q VGND VGND VPWR VPWR final_adder.U$$235/B1 final_adder.U$$729/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$118 _542_/Q _414_/Q VGND VGND VPWR VPWR final_adder.U$$613/B1 final_adder.U$$740/A
+ sky130_fd_sc_hd__ha_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$129 final_adder.U$$623/A final_adder.U$$623/B final_adder.U$$129/B1
+ VGND VGND VPWR VPWR final_adder.U$$624/B sky130_fd_sc_hd__a21o_2
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater388 U$$826/X VGND VGND VPWR VPWR U$$928/A2 sky130_fd_sc_hd__buf_12
XU$$4070 U$$4070/A U$$4109/A VGND VGND VPWR VPWR U$$4070/X sky130_fd_sc_hd__xor2_1
XU$$4081 U$$4492/A1 U$$4107/A2 U$$4494/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4082/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater399 U$$4045/A2 VGND VGND VPWR VPWR U$$4107/A2 sky130_fd_sc_hd__buf_12
XU$$4092 U$$4092/A U$$4109/A VGND VGND VPWR VPWR U$$4092/X sky130_fd_sc_hd__xor2_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3380 _594_/Q U$$3292/X _595_/Q U$$3293/X VGND VGND VPWR VPWR U$$3381/A sky130_fd_sc_hd__a22o_1
XFILLER_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3391 U$$3391/A U$$3403/B VGND VGND VPWR VPWR U$$3391/X sky130_fd_sc_hd__xor2_1
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2690 U$$2690/A _655_/Q VGND VGND VPWR VPWR U$$2690/X sky130_fd_sc_hd__xor2_1
XFILLER_90_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_81_1 dadda_fa_4_81_1/A dadda_fa_4_81_1/B dadda_fa_4_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/B dadda_fa_5_81_1/B sky130_fd_sc_hd__fa_2
Xdadda_fa_4_74_0 dadda_fa_4_74_0/A dadda_fa_4_74_0/B dadda_fa_4_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/A dadda_fa_5_74_1/A sky130_fd_sc_hd__fa_1
XFILLER_1_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput103 b[44] VGND VGND VPWR VPWR _596_/D sky130_fd_sc_hd__clkbuf_1
Xinput114 b[54] VGND VGND VPWR VPWR _606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput125 b[6] VGND VGND VPWR VPWR _558_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput136 c[106] VGND VGND VPWR VPWR input136/X sky130_fd_sc_hd__clkbuf_1
Xinput147 c[116] VGND VGND VPWR VPWR input147/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput158 c[126] VGND VGND VPWR VPWR input158/X sky130_fd_sc_hd__buf_2
Xinput169 c[20] VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$630 final_adder.U$$8/SUM final_adder.U$$630/B VGND VGND VPWR VPWR
+ hold6/A sky130_fd_sc_hd__xor2_2
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$641 final_adder.U$$641/A final_adder.U$$641/B VGND VGND VPWR VPWR
+ _187_/D sky130_fd_sc_hd__xor2_1
X_641_ _679_/CLK _641_/D VGND VGND VPWR VPWR _641_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$652 final_adder.U$$652/A final_adder.U$$652/B VGND VGND VPWR VPWR
+ _198_/D sky130_fd_sc_hd__xor2_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_808__860 VGND VGND VPWR VPWR _808__860/HI U$$4461/B sky130_fd_sc_hd__conb_1
XFILLER_57_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$663 final_adder.U$$663/A final_adder.U$$663/B VGND VGND VPWR VPWR
+ hold5/A sky130_fd_sc_hd__xor2_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$502 U$$502/A U$$547/A VGND VGND VPWR VPWR U$$502/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$674 final_adder.U$$674/A final_adder.U$$674/B VGND VGND VPWR VPWR
+ _220_/D sky130_fd_sc_hd__xor2_1
XFILLER_186_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$513 U$$924/A1 U$$545/A2 U$$926/A1 U$$416/X VGND VGND VPWR VPWR U$$514/A sky130_fd_sc_hd__a22o_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$685 final_adder.U$$685/A final_adder.U$$685/B VGND VGND VPWR VPWR
+ _231_/D sky130_fd_sc_hd__xor2_1
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$524 U$$524/A U$$530/B VGND VGND VPWR VPWR U$$524/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$696 final_adder.U$$696/A final_adder.U$$696/B VGND VGND VPWR VPWR
+ _242_/D sky130_fd_sc_hd__xor2_1
XFILLER_186_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$535 U$$946/A1 U$$415/X U$$948/A1 U$$416/X VGND VGND VPWR VPWR U$$536/A sky130_fd_sc_hd__a22o_1
X_572_ _645_/CLK _572_/D VGND VGND VPWR VPWR _572_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$546 U$$546/A U$$547/A VGND VGND VPWR VPWR U$$546/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$557 U$$557/A U$$623/B VGND VGND VPWR VPWR U$$557/X sky130_fd_sc_hd__xor2_1
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$568 U$$842/A1 U$$626/A2 U$$22/A1 U$$553/X VGND VGND VPWR VPWR U$$569/A sky130_fd_sc_hd__a22o_1
XU$$579 U$$579/A U$$623/B VGND VGND VPWR VPWR U$$579/X sky130_fd_sc_hd__xor2_1
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_89_0 dadda_fa_6_89_0/A dadda_fa_6_89_0/B dadda_fa_6_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_90_0/B dadda_fa_7_89_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_158_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1230 U$$819/A1 U$$1100/X U$$1230/B1 U$$1101/X VGND VGND VPWR VPWR U$$1231/A sky130_fd_sc_hd__a22o_1
XFILLER_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1241 _552_/Q U$$1237/X U$$969/A1 U$$1238/X VGND VGND VPWR VPWR U$$1242/A sky130_fd_sc_hd__a22o_1
XU$$1252 U$$1252/A U$$1336/B VGND VGND VPWR VPWR U$$1252/X sky130_fd_sc_hd__xor2_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1263 U$$28/B1 U$$1237/X U$$32/A1 U$$1238/X VGND VGND VPWR VPWR U$$1264/A sky130_fd_sc_hd__a22o_1
XU$$1274 U$$1274/A U$$1342/B VGND VGND VPWR VPWR U$$1274/X sky130_fd_sc_hd__xor2_1
XFILLER_31_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1285 U$$50/B1 U$$1341/A2 U$$876/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1286/A sky130_fd_sc_hd__a22o_1
XU$$1296 U$$1296/A U$$1342/B VGND VGND VPWR VPWR U$$1296/X sky130_fd_sc_hd__xor2_1
XFILLER_188_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_91_0 dadda_fa_5_91_0/A dadda_fa_5_91_0/B dadda_fa_5_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/A dadda_fa_6_91_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_76_6 U$$3883/X U$$4016/X U$$4149/X VGND VGND VPWR VPWR dadda_fa_2_77_2/B
+ dadda_fa_2_76_5/B sky130_fd_sc_hd__fa_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_69_5 U$$4401/X input222/X dadda_fa_1_69_5/CIN VGND VGND VPWR VPWR dadda_fa_2_70_2/A
+ dadda_fa_2_69_5/A sky130_fd_sc_hd__fa_2
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_96_0 _705__925/HI U$$2327/X VGND VGND VPWR VPWR dadda_fa_3_97_0/A dadda_fa_3_96_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_100_1 dadda_fa_3_100_1/A dadda_fa_3_100_1/B dadda_fa_3_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_0/CIN dadda_fa_4_100_2/A sky130_fd_sc_hd__fa_1
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_121_0 dadda_fa_6_121_0/A dadda_fa_6_121_0/B dadda_fa_6_121_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_122_0/B dadda_fa_7_121_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_64_4 U$$1731/X U$$1864/X U$$1997/X VGND VGND VPWR VPWR dadda_fa_1_65_6/CIN
+ dadda_fa_1_64_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_41_3 dadda_fa_3_41_3/A dadda_fa_3_41_3/B dadda_fa_3_41_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/B dadda_fa_4_41_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$471 final_adder.U$$294/B final_adder.U$$698/B final_adder.U$$205/X
+ VGND VGND VPWR VPWR final_adder.U$$700/B sky130_fd_sc_hd__a21o_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$310 U$$36/A1 U$$278/X U$$38/A1 U$$279/X VGND VGND VPWR VPWR U$$311/A sky130_fd_sc_hd__a22o_1
XFILLER_57_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ _644_/CLK _624_/D VGND VGND VPWR VPWR _624_/Q sky130_fd_sc_hd__dfxtp_4
XU$$321 U$$321/A U$$391/B VGND VGND VPWR VPWR U$$321/X sky130_fd_sc_hd__xor2_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_34_2 dadda_fa_3_34_2/A dadda_fa_3_34_2/B dadda_fa_3_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/A dadda_fa_4_34_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$493 final_adder.U$$316/B final_adder.U$$742/B final_adder.U$$249/X
+ VGND VGND VPWR VPWR final_adder.U$$744/B sky130_fd_sc_hd__a21o_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$332 U$$58/A1 U$$278/X U$$60/A1 U$$279/X VGND VGND VPWR VPWR U$$333/A sky130_fd_sc_hd__a22o_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$343 U$$343/A U$$357/B VGND VGND VPWR VPWR U$$343/X sky130_fd_sc_hd__xor2_2
XFILLER_189_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$354 U$$80/A1 U$$278/X U$$82/A1 U$$279/X VGND VGND VPWR VPWR U$$355/A sky130_fd_sc_hd__a22o_1
XFILLER_189_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$365 U$$365/A U$$391/B VGND VGND VPWR VPWR U$$365/X sky130_fd_sc_hd__xor2_1
XFILLER_17_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_27_1 U$$1524/X U$$1657/X U$$1790/X VGND VGND VPWR VPWR dadda_fa_4_28_0/CIN
+ dadda_fa_4_27_2/A sky130_fd_sc_hd__fa_2
X_555_ _578_/CLK _555_/D VGND VGND VPWR VPWR _555_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$376 U$$924/A1 U$$278/X U$$926/A1 U$$279/X VGND VGND VPWR VPWR U$$377/A sky130_fd_sc_hd__a22o_1
XFILLER_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$387 U$$387/A _621_/Q VGND VGND VPWR VPWR U$$387/X sky130_fd_sc_hd__xor2_2
XU$$398 U$$946/A1 U$$278/X U$$948/A1 U$$279/X VGND VGND VPWR VPWR U$$399/A sky130_fd_sc_hd__a22o_1
XFILLER_60_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_486_ _490_/CLK _486_/D VGND VGND VPWR VPWR _486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_86_5 dadda_fa_2_86_5/A dadda_fa_2_86_5/B dadda_fa_2_86_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_2/A dadda_fa_4_86_0/A sky130_fd_sc_hd__fa_2
XFILLER_153_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_79_4 dadda_fa_2_79_4/A dadda_fa_2_79_4/B dadda_fa_2_79_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/CIN dadda_fa_3_79_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1060 U$$1060/A _631_/Q VGND VGND VPWR VPWR U$$1060/X sky130_fd_sc_hd__xor2_1
XU$$1071 U$$934/A1 U$$963/X U$$799/A1 U$$964/X VGND VGND VPWR VPWR U$$1072/A sky130_fd_sc_hd__a22o_1
XFILLER_148_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1082 U$$1082/A _631_/Q VGND VGND VPWR VPWR U$$1082/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1093 _615_/Q U$$1093/A2 U$$1093/B1 U$$964/X VGND VGND VPWR VPWR U$$1094/A sky130_fd_sc_hd__a22o_1
XFILLER_32_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_116_1 dadda_fa_5_116_1/A dadda_fa_5_116_1/B dadda_fa_5_116_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/B dadda_fa_7_116_0/A sky130_fd_sc_hd__fa_2
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_109_0 dadda_fa_5_109_0/A dadda_fa_5_109_0/B dadda_fa_5_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/A dadda_fa_6_109_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_4 U$$2829/X U$$2962/X U$$3095/X VGND VGND VPWR VPWR dadda_fa_2_82_2/B
+ dadda_fa_2_81_5/A sky130_fd_sc_hd__fa_2
XFILLER_105_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_74_3 U$$2948/X U$$3081/X U$$3214/X VGND VGND VPWR VPWR dadda_fa_2_75_1/B
+ dadda_fa_2_74_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_51_2 dadda_fa_4_51_2/A dadda_fa_4_51_2/B dadda_fa_4_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/CIN dadda_fa_5_51_1/CIN sky130_fd_sc_hd__fa_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_2 U$$3333/X U$$3466/X U$$3599/X VGND VGND VPWR VPWR dadda_fa_2_68_1/A
+ dadda_fa_2_67_4/A sky130_fd_sc_hd__fa_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_1 dadda_fa_4_44_1/A dadda_fa_4_44_1/B dadda_fa_4_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/B dadda_fa_5_44_1/B sky130_fd_sc_hd__fa_1
XFILLER_101_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_21_0 dadda_fa_7_21_0/A dadda_fa_7_21_0/B dadda_fa_7_21_0/CIN VGND VGND
+ VPWR VPWR _446_/D _317_/D sky130_fd_sc_hd__fa_2
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_37_0 dadda_fa_4_37_0/A dadda_fa_4_37_0/B dadda_fa_4_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/A dadda_fa_5_37_1/A sky130_fd_sc_hd__fa_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _480_/CLK _340_/D VGND VGND VPWR VPWR _340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_271_ _280_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_0_70_4 U$$2009/X U$$2142/X VGND VGND VPWR VPWR dadda_fa_1_71_7/CIN dadda_fa_2_70_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_185_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_89_3 dadda_fa_3_89_3/A dadda_fa_3_89_3/B dadda_fa_3_89_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/B dadda_fa_4_89_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_2_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_56_2 U$$917/X U$$1050/X VGND VGND VPWR VPWR dadda_fa_1_57_8/A dadda_fa_2_56_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_1_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_62_1 U$$530/X U$$663/X U$$796/X VGND VGND VPWR VPWR dadda_fa_1_63_5/CIN
+ dadda_fa_1_62_7/CIN sky130_fd_sc_hd__fa_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3902 _581_/Q U$$3912/A2 _582_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3903/A sky130_fd_sc_hd__a22o_1
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_55_0 U$$117/X U$$250/X U$$383/X VGND VGND VPWR VPWR dadda_fa_1_56_7/CIN
+ dadda_fa_1_55_8/CIN sky130_fd_sc_hd__fa_2
XU$$3913 U$$3913/A U$$3929/B VGND VGND VPWR VPWR U$$3913/X sky130_fd_sc_hd__xor2_1
XU$$3924 U$$4335/A1 U$$3840/X _593_/Q U$$3841/X VGND VGND VPWR VPWR U$$3925/A sky130_fd_sc_hd__a22o_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3935 U$$3935/A _673_/Q VGND VGND VPWR VPWR U$$3935/X sky130_fd_sc_hd__xor2_1
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3946 U$$4494/A1 U$$3970/A2 U$$4496/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3947/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3957 U$$3957/A _673_/Q VGND VGND VPWR VPWR U$$3957/X sky130_fd_sc_hd__xor2_1
XFILLER_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$290 final_adder.U$$290/A final_adder.U$$290/B VGND VGND VPWR VPWR
+ final_adder.U$$336/A sky130_fd_sc_hd__and2_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$140 U$$274/A U$$140/B VGND VGND VPWR VPWR U$$140/X sky130_fd_sc_hd__and2_1
XU$$3968 U$$4379/A1 U$$3970/A2 U$$819/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3969/A
+ sky130_fd_sc_hd__a22o_1
X_607_ _611_/CLK _607_/D VGND VGND VPWR VPWR _607_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$151 U$$12/B1 U$$141/X U$$16/A1 U$$142/X VGND VGND VPWR VPWR U$$152/A sky130_fd_sc_hd__a22o_1
XU$$3979 U$$3979/A1 U$$3977/X U$$4255/A1 U$$3978/X VGND VGND VPWR VPWR U$$3980/A sky130_fd_sc_hd__a22o_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$162 U$$162/A U$$274/A VGND VGND VPWR VPWR U$$162/X sky130_fd_sc_hd__xor2_1
XU$$173 U$$36/A1 U$$141/X U$$38/A1 U$$142/X VGND VGND VPWR VPWR U$$174/A sky130_fd_sc_hd__a22o_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$184 U$$184/A U$$242/B VGND VGND VPWR VPWR U$$184/X sky130_fd_sc_hd__xor2_1
XFILLER_72_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$195 U$$58/A1 U$$141/X U$$60/A1 U$$142/X VGND VGND VPWR VPWR U$$196/A sky130_fd_sc_hd__a22o_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_538_ _595_/CLK _538_/D VGND VGND VPWR VPWR _538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_469_ _469_/CLK _469_/D VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_91_3 U$$4312/X U$$4445/X input247/X VGND VGND VPWR VPWR dadda_fa_3_92_1/B
+ dadda_fa_3_91_3/B sky130_fd_sc_hd__fa_2
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_84_2 dadda_fa_2_84_2/A dadda_fa_2_84_2/B dadda_fa_2_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/A dadda_fa_3_84_3/A sky130_fd_sc_hd__fa_1
XFILLER_5_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput259 _269_/Q VGND VGND VPWR VPWR o[101] sky130_fd_sc_hd__buf_2
X_713__765 VGND VGND VPWR VPWR _713__765/HI U$$1230/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_5_61_1 dadda_fa_5_61_1/A dadda_fa_5_61_1/B dadda_fa_5_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/B dadda_fa_7_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_77_1 dadda_fa_2_77_1/A dadda_fa_2_77_1/B dadda_fa_2_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/CIN dadda_fa_3_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_54_0 dadda_fa_5_54_0/A dadda_fa_5_54_0/B dadda_fa_5_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/A dadda_fa_6_54_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_53_8 U$$3571/X input205/X dadda_fa_1_53_8/CIN VGND VGND VPWR VPWR dadda_fa_2_54_3/A
+ dadda_fa_3_53_0/A sky130_fd_sc_hd__fa_2
XFILLER_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_100_0 _693__913/HI U$$2601/X U$$2734/X VGND VGND VPWR VPWR dadda_fa_3_101_1/B
+ dadda_fa_3_100_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_99_2 dadda_fa_4_99_2/A dadda_fa_4_99_2/B dadda_fa_4_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/CIN dadda_fa_5_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_69_0 dadda_fa_7_69_0/A dadda_fa_7_69_0/B dadda_fa_7_69_0/CIN VGND VGND
+ VPWR VPWR _494_/D _365_/D sky130_fd_sc_hd__fa_2
XFILLER_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_72_0 U$$2013/X U$$2146/X U$$2279/X VGND VGND VPWR VPWR dadda_fa_2_73_0/B
+ dadda_fa_2_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_87_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3209 U$$4442/A1 U$$3243/A2 U$$4170/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3210/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2508 U$$4289/A1 U$$2534/A2 U$$4289/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2509/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2519 U$$2519/A U$$2585/B VGND VGND VPWR VPWR U$$2519/X sky130_fd_sc_hd__xor2_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1807 U$$4273/A1 U$$1903/A2 U$$987/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1808/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_703__923 VGND VGND VPWR VPWR _703__923/HI _703__923/LO sky130_fd_sc_hd__conb_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1818 U$$1818/A U$$1918/A VGND VGND VPWR VPWR U$$1818/X sky130_fd_sc_hd__xor2_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1829 U$$48/A1 U$$1897/A2 U$$50/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1830/A sky130_fd_sc_hd__a22o_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_323_ _333_/CLK _323_/D VGND VGND VPWR VPWR _323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254_ _503_/CLK _254_/D VGND VGND VPWR VPWR _254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_185_ _333_/CLK _185_/D VGND VGND VPWR VPWR _185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_94_1 dadda_fa_3_94_1/A dadda_fa_3_94_1/B dadda_fa_3_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/CIN dadda_fa_4_94_2/A sky130_fd_sc_hd__fa_2
XFILLER_171_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_71_0 dadda_fa_6_71_0/A dadda_fa_6_71_0/B dadda_fa_6_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_72_0/B dadda_fa_7_71_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_170_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_87_0 dadda_fa_3_87_0/A dadda_fa_3_87_0/B dadda_fa_3_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/B dadda_fa_4_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater707 U$$54/A1 VGND VGND VPWR VPWR U$$876/A1 sky130_fd_sc_hd__buf_12
XU$$4400 _556_/Q U$$4388/X _557_/Q U$$4389/X VGND VGND VPWR VPWR U$$4401/A sky130_fd_sc_hd__a22o_1
Xrepeater718 U$$46/A1 VGND VGND VPWR VPWR U$$4291/B1 sky130_fd_sc_hd__buf_12
XU$$4411 U$$4411/A U$$4411/B VGND VGND VPWR VPWR U$$4411/X sky130_fd_sc_hd__xor2_1
Xrepeater729 _566_/Q VGND VGND VPWR VPWR U$$4283/A1 sky130_fd_sc_hd__buf_12
XU$$4422 _567_/Q U$$4388/X U$$4424/A1 U$$4389/X VGND VGND VPWR VPWR U$$4423/A sky130_fd_sc_hd__a22o_2
XU$$4433 U$$4433/A U$$4433/B VGND VGND VPWR VPWR U$$4433/X sky130_fd_sc_hd__xor2_1
XU$$4444 _578_/Q U$$4388/X U$$4446/A1 U$$4389/X VGND VGND VPWR VPWR U$$4445/A sky130_fd_sc_hd__a22o_1
XU$$3710 U$$3710/A U$$3784/B VGND VGND VPWR VPWR U$$3710/X sky130_fd_sc_hd__xor2_1
XU$$4455 U$$4455/A U$$4455/B VGND VGND VPWR VPWR U$$4455/X sky130_fd_sc_hd__xor2_2
XU$$3721 U$$22/A1 U$$3795/A2 U$$4271/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3722/A sky130_fd_sc_hd__a22o_1
XU$$4466 U$$82/A1 U$$4388/X U$$632/A1 U$$4389/X VGND VGND VPWR VPWR U$$4467/A sky130_fd_sc_hd__a22o_2
Xdadda_fa_4_116_0 U$$3830/X U$$3963/X U$$4096/X VGND VGND VPWR VPWR dadda_fa_5_117_0/A
+ dadda_fa_5_116_1/A sky130_fd_sc_hd__fa_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_49_5 dadda_fa_2_49_5/A dadda_fa_2_49_5/B dadda_fa_2_49_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_2/A dadda_fa_4_49_0/A sky130_fd_sc_hd__fa_2
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4477 U$$4477/A U$$4477/B VGND VGND VPWR VPWR U$$4477/X sky130_fd_sc_hd__xor2_1
XFILLER_93_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3732 U$$3732/A U$$3756/B VGND VGND VPWR VPWR U$$3732/X sky130_fd_sc_hd__xor2_1
XU$$3743 U$$4289/B1 U$$3795/A2 U$$4291/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3744/A
+ sky130_fd_sc_hd__a22o_1
XU$$4488 U$$787/B1 U$$4388/X U$$654/A1 U$$4389/X VGND VGND VPWR VPWR U$$4489/A sky130_fd_sc_hd__a22o_1
XFILLER_65_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3754 U$$3754/A U$$3794/B VGND VGND VPWR VPWR U$$3754/X sky130_fd_sc_hd__xor2_1
XU$$4499 U$$4499/A U$$4499/B VGND VGND VPWR VPWR U$$4499/X sky130_fd_sc_hd__xor2_2
XU$$3765 _581_/Q U$$3783/A2 _582_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3766/A sky130_fd_sc_hd__a22o_1
XU$$3776 U$$3776/A U$$3794/B VGND VGND VPWR VPWR U$$3776/X sky130_fd_sc_hd__xor2_2
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3787 U$$4335/A1 U$$3795/A2 _593_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3788/A sky130_fd_sc_hd__a22o_1
XFILLER_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3798 U$$3798/A _671_/Q VGND VGND VPWR VPWR U$$3798/X sky130_fd_sc_hd__xor2_1
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_51_5 U$$2104/X U$$2237/X U$$2370/X VGND VGND VPWR VPWR dadda_fa_2_52_2/A
+ dadda_fa_2_51_5/A sky130_fd_sc_hd__fa_2
XFILLER_68_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$909 U$$909/A U$$943/B VGND VGND VPWR VPWR U$$909/X sky130_fd_sc_hd__xor2_1
XFILLER_141_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_44_4 U$$1691/X U$$1824/X U$$1957/X VGND VGND VPWR VPWR dadda_fa_2_45_3/CIN
+ dadda_fa_2_44_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_55_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_841__893 VGND VGND VPWR VPWR _841__893/HI U$$682/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_14_2 U$$998/B input162/X dadda_ha_3_14_0/SUM VGND VGND VPWR VPWR dadda_fa_5_15_0/CIN
+ dadda_fa_5_14_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_19_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3006 U$$3006/A _659_/Q VGND VGND VPWR VPWR U$$3006/X sky130_fd_sc_hd__xor2_1
XFILLER_189_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3017 _661_/Q U$$3017/B VGND VGND VPWR VPWR U$$3017/X sky130_fd_sc_hd__and2_1
XFILLER_35_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3028 _555_/Q U$$3146/A2 _556_/Q U$$3146/B2 VGND VGND VPWR VPWR U$$3029/A sky130_fd_sc_hd__a22o_1
XU$$3039 U$$3039/A U$$3085/B VGND VGND VPWR VPWR U$$3039/X sky130_fd_sc_hd__xor2_1
XFILLER_35_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2305 U$$2305/A U$$2327/B VGND VGND VPWR VPWR U$$2305/X sky130_fd_sc_hd__xor2_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2316 U$$4508/A1 U$$2316/A2 U$$4510/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2317/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2327 U$$2327/A U$$2327/B VGND VGND VPWR VPWR U$$2327/X sky130_fd_sc_hd__xor2_2
XU$$2338 U$$2338/A U$$2432/B VGND VGND VPWR VPWR U$$2338/X sky130_fd_sc_hd__xor2_2
XU$$2349 U$$20/A1 U$$2333/X U$$979/B1 U$$2334/X VGND VGND VPWR VPWR U$$2350/A sky130_fd_sc_hd__a22o_1
XU$$1604 U$$1604/A U$$1614/B VGND VGND VPWR VPWR U$$1604/X sky130_fd_sc_hd__xor2_2
XU$$1615 _602_/Q U$$1641/A2 _603_/Q U$$1641/B2 VGND VGND VPWR VPWR U$$1616/A sky130_fd_sc_hd__a22o_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1626 U$$1626/A U$$1643/A VGND VGND VPWR VPWR U$$1626/X sky130_fd_sc_hd__xor2_1
XU$$1637 _613_/Q U$$1641/A2 _614_/Q U$$1641/B2 VGND VGND VPWR VPWR U$$1638/A sky130_fd_sc_hd__a22o_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1648 U$$1646/Y _640_/Q _639_/Q U$$1647/X U$$1644/Y VGND VGND VPWR VPWR U$$1648/X
+ sky130_fd_sc_hd__a32o_4
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1659 U$$1659/A U$$1781/A VGND VGND VPWR VPWR U$$1659/X sky130_fd_sc_hd__xor2_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ _327_/CLK _306_/D VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_237_ _499_/CLK _237_/D VGND VGND VPWR VPWR _237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_168_ _448_/CLK _168_/D VGND VGND VPWR VPWR _168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_784__836 VGND VGND VPWR VPWR _784__836/HI U$$4413/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_61_4 dadda_fa_2_61_4/A dadda_fa_2_61_4/B dadda_fa_2_61_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/CIN dadda_fa_3_61_3/CIN sky130_fd_sc_hd__fa_2
Xrepeater504 U$$1770/B2 VGND VGND VPWR VPWR U$$1734/B2 sky130_fd_sc_hd__buf_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater515 _679_/Q VGND VGND VPWR VPWR U$$4384/A sky130_fd_sc_hd__buf_12
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater526 U$$3784/B VGND VGND VPWR VPWR U$$3756/B sky130_fd_sc_hd__buf_12
XFILLER_133_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater537 U$$3403/B VGND VGND VPWR VPWR U$$3397/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_54_3 dadda_fa_2_54_3/A dadda_fa_2_54_3/B dadda_fa_2_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/B dadda_fa_3_54_3/B sky130_fd_sc_hd__fa_2
XU$$4230 U$$4504/A1 U$$4244/A2 U$$4506/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4231/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater548 _659_/Q VGND VGND VPWR VPWR U$$3004/B sky130_fd_sc_hd__buf_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater559 _651_/Q VGND VGND VPWR VPWR U$$2436/B sky130_fd_sc_hd__buf_12
XU$$4241 U$$4241/A U$$4246/A VGND VGND VPWR VPWR U$$4241/X sky130_fd_sc_hd__xor2_1
XU$$4252 U$$4250/B U$$4247/A _678_/Q U$$4247/Y VGND VGND VPWR VPWR U$$4252/X sky130_fd_sc_hd__a22o_4
XU$$4263 _556_/Q U$$4381/A2 _557_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4264/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_2 dadda_fa_2_47_2/A dadda_fa_2_47_2/B dadda_fa_2_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/A dadda_fa_3_47_3/A sky130_fd_sc_hd__fa_1
X_825__877 VGND VGND VPWR VPWR _825__877/HI U$$4495/B sky130_fd_sc_hd__conb_1
XU$$4274 U$$4274/A U$$4332/B VGND VGND VPWR VPWR U$$4274/X sky130_fd_sc_hd__xor2_1
XU$$4285 U$$4285/A1 U$$4251/X U$$4424/A1 U$$4252/X VGND VGND VPWR VPWR U$$4286/A sky130_fd_sc_hd__a22o_1
XU$$3540 U$$3540/A U$$3561/A VGND VGND VPWR VPWR U$$3540/X sky130_fd_sc_hd__xor2_1
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3551 U$$4510/A1 U$$3429/X U$$539/A1 U$$3430/X VGND VGND VPWR VPWR U$$3552/A sky130_fd_sc_hd__a22o_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_24_1 dadda_fa_5_24_1/A dadda_fa_5_24_1/B dadda_fa_5_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/B dadda_fa_7_24_0/A sky130_fd_sc_hd__fa_2
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4296 U$$4296/A _679_/Q VGND VGND VPWR VPWR U$$4296/X sky130_fd_sc_hd__xor2_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3562 _667_/Q VGND VGND VPWR VPWR U$$3562/Y sky130_fd_sc_hd__inv_1
XU$$3573 U$$3573/A U$$3625/B VGND VGND VPWR VPWR U$$3573/X sky130_fd_sc_hd__xor2_2
XFILLER_111_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_17_0 dadda_fa_5_17_0/A dadda_fa_5_17_0/B dadda_fa_5_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/A dadda_fa_6_17_0/CIN sky130_fd_sc_hd__fa_1
XU$$3584 U$$22/A1 U$$3624/A2 U$$4271/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3585/A sky130_fd_sc_hd__a22o_1
XU$$2850 _603_/Q U$$2870/A2 _604_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2851/A sky130_fd_sc_hd__a22o_1
XU$$3595 U$$3595/A _669_/Q VGND VGND VPWR VPWR U$$3595/X sky130_fd_sc_hd__xor2_1
XU$$2861 U$$2861/A _657_/Q VGND VGND VPWR VPWR U$$2861/X sky130_fd_sc_hd__xor2_1
XU$$2872 U$$4379/A1 U$$2744/X U$$956/A1 U$$2745/X VGND VGND VPWR VPWR U$$2873/A sky130_fd_sc_hd__a22o_1
XU$$2883 U$$2883/A1 U$$3009/A2 U$$8/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2884/A sky130_fd_sc_hd__a22o_1
XFILLER_178_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2894 U$$2894/A U$$2996/B VGND VGND VPWR VPWR U$$2894/X sky130_fd_sc_hd__xor2_1
XFILLER_179_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_719__771 VGND VGND VPWR VPWR _719__771/HI U$$1504/B1 sky130_fd_sc_hd__conb_1
XFILLER_119_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$706 U$$706/A U$$784/B VGND VGND VPWR VPWR U$$706/X sky130_fd_sc_hd__xor2_2
XU$$717 U$$32/A1 U$$817/A2 U$$34/A1 U$$785/B2 VGND VGND VPWR VPWR U$$718/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_42_1 U$$490/X U$$623/X U$$756/X VGND VGND VPWR VPWR dadda_fa_2_43_3/B
+ dadda_fa_2_42_5/A sky130_fd_sc_hd__fa_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$728 U$$728/A U$$784/B VGND VGND VPWR VPWR U$$728/X sky130_fd_sc_hd__xor2_1
XU$$739 U$$876/A1 U$$785/A2 U$$878/A1 U$$785/B2 VGND VGND VPWR VPWR U$$740/A sky130_fd_sc_hd__a22o_1
XFILLER_44_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_71_3 dadda_fa_3_71_3/A dadda_fa_3_71_3/B dadda_fa_3_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/B dadda_fa_4_71_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_64_2 dadda_fa_3_64_2/A dadda_fa_3_64_2/B dadda_fa_3_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/A dadda_fa_4_64_2/B sky130_fd_sc_hd__fa_1
XFILLER_121_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_57_1 dadda_fa_3_57_1/A dadda_fa_3_57_1/B dadda_fa_3_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/CIN dadda_fa_4_57_2/A sky130_fd_sc_hd__fa_1
XFILLER_117_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_34_0 dadda_fa_6_34_0/A dadda_fa_6_34_0/B dadda_fa_6_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_35_0/B dadda_fa_7_34_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_48_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2102 U$$2102/A U$$2118/B VGND VGND VPWR VPWR U$$2102/X sky130_fd_sc_hd__xor2_1
XFILLER_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2113 U$$880/A1 U$$2117/A2 U$$60/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2114/A sky130_fd_sc_hd__a22o_1
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2124 U$$2124/A _647_/Q VGND VGND VPWR VPWR U$$2124/X sky130_fd_sc_hd__xor2_1
XU$$2135 U$$765/A1 U$$2189/A2 U$$82/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2136/A sky130_fd_sc_hd__a22o_1
XFILLER_90_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1401 U$$1401/A U$$1461/B VGND VGND VPWR VPWR U$$1401/X sky130_fd_sc_hd__xor2_1
XU$$2146 U$$2146/A _647_/Q VGND VGND VPWR VPWR U$$2146/X sky130_fd_sc_hd__xor2_1
XU$$2157 _599_/Q U$$2189/A2 _600_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2158/A sky130_fd_sc_hd__a22o_1
XFILLER_34_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1412 U$$3876/B1 U$$1472/A2 U$$4291/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1413/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2168 U$$2168/A U$$2192/A VGND VGND VPWR VPWR U$$2168/X sky130_fd_sc_hd__xor2_1
XU$$1423 U$$1423/A U$$1461/B VGND VGND VPWR VPWR U$$1423/X sky130_fd_sc_hd__xor2_1
XU$$1434 U$$64/A1 U$$1472/A2 U$$66/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1435/A sky130_fd_sc_hd__a22o_1
XU$$2179 U$$4508/A1 U$$2189/A2 U$$4510/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2180/A
+ sky130_fd_sc_hd__a22o_1
XU$$1445 U$$1445/A U$$1505/B VGND VGND VPWR VPWR U$$1445/X sky130_fd_sc_hd__xor2_1
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1456 U$$86/A1 U$$1472/A2 U$$88/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1457/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1467 U$$1467/A U$$1479/B VGND VGND VPWR VPWR U$$1467/X sky130_fd_sc_hd__xor2_1
XFILLER_43_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1478 U$$930/A1 U$$1374/X U$$932/A1 U$$1375/X VGND VGND VPWR VPWR U$$1479/A sky130_fd_sc_hd__a22o_1
XFILLER_187_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1489 U$$1489/A _637_/Q VGND VGND VPWR VPWR U$$1489/X sky130_fd_sc_hd__xor2_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_107_0 dadda_fa_7_107_0/A dadda_fa_7_107_0/B dadda_fa_7_107_0/CIN VGND
+ VGND VPWR VPWR _532_/D _403_/D sky130_fd_sc_hd__fa_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$108 _532_/Q _404_/Q VGND VGND VPWR VPWR final_adder.U$$603/B1 final_adder.U$$730/A
+ sky130_fd_sc_hd__ha_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$119 _543_/Q _415_/Q VGND VGND VPWR VPWR final_adder.U$$247/B1 final_adder.U$$741/A
+ sky130_fd_sc_hd__ha_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_52_0 dadda_fa_2_52_0/A dadda_fa_2_52_0/B dadda_fa_2_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/B dadda_fa_3_52_2/B sky130_fd_sc_hd__fa_2
XFILLER_111_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater389 U$$817/A2 VGND VGND VPWR VPWR U$$785/A2 sky130_fd_sc_hd__buf_12
XU$$4060 U$$4060/A _675_/Q VGND VGND VPWR VPWR U$$4060/X sky130_fd_sc_hd__xor2_1
XU$$4071 U$$98/A1 U$$4107/A2 U$$4484/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4072/A sky130_fd_sc_hd__a22o_1
XU$$4082 U$$4082/A U$$4109/A VGND VGND VPWR VPWR U$$4082/X sky130_fd_sc_hd__xor2_1
XFILLER_54_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4093 U$$4504/A1 U$$4107/A2 U$$4506/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4094/A
+ sky130_fd_sc_hd__a22o_1
XU$$3370 U$$630/A1 U$$3412/A2 U$$632/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3371/A sky130_fd_sc_hd__a22o_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3381 U$$3381/A U$$3403/B VGND VGND VPWR VPWR U$$3381/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3392 _600_/Q U$$3396/A2 _601_/Q U$$3396/B2 VGND VGND VPWR VPWR U$$3393/A sky130_fd_sc_hd__a22o_1
XU$$2680 U$$2680/A U$$2698/B VGND VGND VPWR VPWR U$$2680/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_6_0 U$$19/X U$$152/X U$$285/X VGND VGND VPWR VPWR dadda_fa_6_7_0/A dadda_fa_6_6_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_178_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2691 U$$771/B1 U$$2729/A2 U$$912/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2692/A sky130_fd_sc_hd__a22o_1
XFILLER_90_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_60_clk _536_/CLK VGND VGND VPWR VPWR _614_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1990 U$$892/B1 U$$2036/A2 U$$74/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1991/A sky130_fd_sc_hd__a22o_1
XFILLER_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_81_2 dadda_fa_4_81_2/A dadda_fa_4_81_2/B dadda_fa_4_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/CIN dadda_fa_5_81_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_74_1 dadda_fa_4_74_1/A dadda_fa_4_74_1/B dadda_fa_4_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/B dadda_fa_5_74_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_51_0 dadda_fa_7_51_0/A dadda_fa_7_51_0/B dadda_fa_7_51_0/CIN VGND VGND
+ VPWR VPWR _476_/D _347_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_67_0 dadda_fa_4_67_0/A dadda_fa_4_67_0/B dadda_fa_4_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/A dadda_fa_5_67_1/A sky130_fd_sc_hd__fa_1
Xinput104 b[45] VGND VGND VPWR VPWR _597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput115 b[55] VGND VGND VPWR VPWR _607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput126 b[7] VGND VGND VPWR VPWR _559_/D sky130_fd_sc_hd__buf_4
Xinput137 c[107] VGND VGND VPWR VPWR input137/X sky130_fd_sc_hd__buf_2
Xinput148 c[117] VGND VGND VPWR VPWR input148/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput159 c[127] VGND VGND VPWR VPWR input159/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$631 final_adder.U$$9/SUM final_adder.U$$631/B VGND VGND VPWR VPWR
+ _177_/D sky130_fd_sc_hd__xor2_2
X_640_ _647_/CLK _640_/D VGND VGND VPWR VPWR _640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$642 final_adder.U$$642/A final_adder.U$$642/B VGND VGND VPWR VPWR
+ _188_/D sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$653 final_adder.U$$653/A final_adder.U$$653/B VGND VGND VPWR VPWR
+ _199_/D sky130_fd_sc_hd__xor2_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$664 final_adder.U$$664/A final_adder.U$$664/B VGND VGND VPWR VPWR
+ _210_/D sky130_fd_sc_hd__xor2_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$503 U$$92/A1 U$$545/A2 U$$92/B1 U$$416/X VGND VGND VPWR VPWR U$$504/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$675 final_adder.U$$675/A final_adder.U$$675/B VGND VGND VPWR VPWR
+ _221_/D sky130_fd_sc_hd__xor2_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$514 U$$514/A U$$547/A VGND VGND VPWR VPWR U$$514/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$686 final_adder.U$$686/A final_adder.U$$686/B VGND VGND VPWR VPWR
+ hold2/A sky130_fd_sc_hd__xor2_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$525 U$$799/A1 U$$545/A2 U$$938/A1 U$$416/X VGND VGND VPWR VPWR U$$526/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_571_ _576_/CLK _571_/D VGND VGND VPWR VPWR _571_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$697 final_adder.U$$697/A final_adder.U$$697/B VGND VGND VPWR VPWR
+ _243_/D sky130_fd_sc_hd__xor2_1
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$536 U$$536/A _623_/Q VGND VGND VPWR VPWR U$$536/X sky130_fd_sc_hd__xor2_1
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$547 U$$547/A VGND VGND VPWR VPWR U$$547/Y sky130_fd_sc_hd__inv_1
XFILLER_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$558 U$$969/A1 U$$626/A2 U$$971/A1 U$$553/X VGND VGND VPWR VPWR U$$559/A sky130_fd_sc_hd__a22o_1
XU$$569 U$$569/A U$$623/B VGND VGND VPWR VPWR U$$569/X sky130_fd_sc_hd__xor2_1
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk _536_/CLK VGND VGND VPWR VPWR _615_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1220 _610_/Q U$$1100/X U$$4510/A1 U$$1101/X VGND VGND VPWR VPWR U$$1221/A sky130_fd_sc_hd__a22o_1
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1231 U$$1231/A _633_/Q VGND VGND VPWR VPWR U$$1231/X sky130_fd_sc_hd__xor2_1
XU$$1242 U$$1242/A U$$1336/B VGND VGND VPWR VPWR U$$1242/X sky130_fd_sc_hd__xor2_1
XU$$1253 U$$20/A1 U$$1237/X _559_/Q U$$1238/X VGND VGND VPWR VPWR U$$1254/A sky130_fd_sc_hd__a22o_1
XU$$1264 U$$1264/A U$$1336/B VGND VGND VPWR VPWR U$$1264/X sky130_fd_sc_hd__xor2_1
XFILLER_188_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _387_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1275 U$$3876/B1 U$$1341/A2 U$$4291/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1276/A
+ sky130_fd_sc_hd__a22o_1
XU$$1286 U$$1286/A U$$1342/B VGND VGND VPWR VPWR U$$1286/X sky130_fd_sc_hd__xor2_1
XU$$1297 U$$64/A1 U$$1341/A2 U$$66/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1298/A sky130_fd_sc_hd__a22o_1
XFILLER_102_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_91_1 dadda_fa_5_91_1/A dadda_fa_5_91_1/B dadda_fa_5_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/B dadda_fa_7_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_102_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_84_0 dadda_fa_5_84_0/A dadda_fa_5_84_0/B dadda_fa_5_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/A dadda_fa_6_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_76_7 U$$4282/X U$$4415/X input230/X VGND VGND VPWR VPWR dadda_fa_2_77_2/CIN
+ dadda_fa_2_76_5/CIN sky130_fd_sc_hd__fa_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_6 dadda_fa_1_69_6/A dadda_fa_1_69_6/B dadda_fa_1_69_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/B dadda_fa_2_69_5/B sky130_fd_sc_hd__fa_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_99_0 dadda_fa_7_99_0/A dadda_fa_7_99_0/B dadda_fa_7_99_0/CIN VGND VGND
+ VPWR VPWR _524_/D _395_/D sky130_fd_sc_hd__fa_2
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_100_2 dadda_fa_3_100_2/A dadda_fa_3_100_2/B dadda_fa_3_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/A dadda_fa_4_100_2/B sky130_fd_sc_hd__fa_1
XFILLER_107_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_64_5 U$$2130/X U$$2263/X U$$2396/X VGND VGND VPWR VPWR dadda_fa_1_65_7/A
+ dadda_fa_2_64_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_6_114_0 dadda_fa_6_114_0/A dadda_fa_6_114_0/B dadda_fa_6_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_115_0/B dadda_fa_7_114_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$300 U$$26/A1 U$$278/X U$$987/A1 U$$279/X VGND VGND VPWR VPWR U$$301/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$461 final_adder.U$$284/B final_adder.U$$678/B final_adder.U$$185/X
+ VGND VGND VPWR VPWR final_adder.U$$680/B sky130_fd_sc_hd__a21o_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_623_ _644_/CLK _623_/D VGND VGND VPWR VPWR _623_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$311 U$$311/A U$$391/B VGND VGND VPWR VPWR U$$311/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$483 final_adder.U$$306/B final_adder.U$$722/B final_adder.U$$229/X
+ VGND VGND VPWR VPWR final_adder.U$$724/B sky130_fd_sc_hd__a21o_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_34_3 dadda_fa_3_34_3/A dadda_fa_3_34_3/B dadda_fa_3_34_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/B dadda_fa_4_34_2/CIN sky130_fd_sc_hd__fa_2
XU$$322 _572_/Q U$$278/X U$$735/A1 U$$279/X VGND VGND VPWR VPWR U$$323/A sky130_fd_sc_hd__a22o_1
XFILLER_57_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$333 U$$333/A U$$391/B VGND VGND VPWR VPWR U$$333/X sky130_fd_sc_hd__xor2_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$344 U$$68/B1 U$$278/X U$$70/B1 U$$279/X VGND VGND VPWR VPWR U$$345/A sky130_fd_sc_hd__a22o_1
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_2 input176/X dadda_fa_3_27_2/B dadda_fa_3_27_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_28_1/A dadda_fa_4_27_2/B sky130_fd_sc_hd__fa_2
XU$$355 U$$355/A _621_/Q VGND VGND VPWR VPWR U$$355/X sky130_fd_sc_hd__xor2_1
XFILLER_33_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_554_ _573_/CLK _554_/D VGND VGND VPWR VPWR _554_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$366 U$$92/A1 U$$278/X U$$94/A1 U$$279/X VGND VGND VPWR VPWR U$$367/A sky130_fd_sc_hd__a22o_1
XFILLER_33_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$377 U$$377/A _621_/Q VGND VGND VPWR VPWR U$$377/X sky130_fd_sc_hd__xor2_2
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$388 U$$799/A1 U$$278/X U$$938/A1 U$$279/X VGND VGND VPWR VPWR U$$389/A sky130_fd_sc_hd__a22o_1
XU$$399 U$$399/A _621_/Q VGND VGND VPWR VPWR U$$399/X sky130_fd_sc_hd__xor2_1
XFILLER_72_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_485_ _490_/CLK _485_/D VGND VGND VPWR VPWR _485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk _369_/CLK VGND VGND VPWR VPWR _476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_79_5 dadda_fa_2_79_5/A dadda_fa_2_79_5/B dadda_fa_2_79_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_2/A dadda_fa_4_79_0/A sky130_fd_sc_hd__fa_2
XFILLER_113_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_2_30_4 U$$1663/X U$$1796/X VGND VGND VPWR VPWR dadda_fa_3_31_2/B dadda_fa_4_30_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_132_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_7_0_0 U$$7/X U$$9/B VGND VGND VPWR VPWR _425_/D _296_/D sky130_fd_sc_hd__ha_2
XFILLER_36_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _464_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1050 U$$1050/A U$$980/B VGND VGND VPWR VPWR U$$1050/X sky130_fd_sc_hd__xor2_1
XU$$1061 U$$924/A1 U$$1093/A2 U$$926/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1062/A sky130_fd_sc_hd__a22o_1
XFILLER_52_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1072 U$$1072/A _631_/Q VGND VGND VPWR VPWR U$$1072/X sky130_fd_sc_hd__xor2_1
XU$$1083 U$$946/A1 U$$963/X U$$948/A1 U$$964/X VGND VGND VPWR VPWR U$$1084/A sky130_fd_sc_hd__a22o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1094 U$$1094/A _631_/Q VGND VGND VPWR VPWR U$$1094/X sky130_fd_sc_hd__xor2_1
XFILLER_188_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_82_7 U$$4028/X U$$4161/X VGND VGND VPWR VPWR dadda_fa_2_83_3/CIN dadda_fa_3_82_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_191_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_109_1 dadda_fa_5_109_1/A dadda_fa_5_109_1/B dadda_fa_5_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/B dadda_fa_7_109_0/A sky130_fd_sc_hd__fa_2
XFILLER_176_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_81_5 U$$3228/X U$$3361/X U$$3494/X VGND VGND VPWR VPWR dadda_fa_2_82_2/CIN
+ dadda_fa_2_81_5/B sky130_fd_sc_hd__fa_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_74_4 U$$3347/X U$$3480/X U$$3613/X VGND VGND VPWR VPWR dadda_fa_2_75_1/CIN
+ dadda_fa_2_74_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_67_3 U$$3732/X U$$3865/X U$$3998/X VGND VGND VPWR VPWR dadda_fa_2_68_1/B
+ dadda_fa_2_67_4/B sky130_fd_sc_hd__fa_1
XFILLER_112_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_2 dadda_fa_4_44_2/A dadda_fa_4_44_2/B dadda_fa_4_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/CIN dadda_fa_5_44_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_1 dadda_fa_4_37_1/A dadda_fa_4_37_1/B dadda_fa_4_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/B dadda_fa_5_37_1/B sky130_fd_sc_hd__fa_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_14_0 dadda_fa_7_14_0/A dadda_fa_7_14_0/B dadda_fa_7_14_0/CIN VGND VGND
+ VPWR VPWR _439_/D _310_/D sky130_fd_sc_hd__fa_2
XFILLER_148_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_270_ _280_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_62_2 U$$929/X U$$1062/X U$$1195/X VGND VGND VPWR VPWR dadda_fa_1_63_6/A
+ dadda_fa_1_62_8/A sky130_fd_sc_hd__fa_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3903 U$$3903/A U$$3929/B VGND VGND VPWR VPWR U$$3903/X sky130_fd_sc_hd__xor2_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3914 U$$78/A1 U$$3970/A2 U$$765/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3915/A sky130_fd_sc_hd__a22o_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3925 U$$3925/A U$$3929/B VGND VGND VPWR VPWR U$$3925/X sky130_fd_sc_hd__xor2_1
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3936 U$$4484/A1 U$$3970/A2 U$$4486/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3937/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_32_0 U$$2289/B input182/X dadda_fa_3_32_0/CIN VGND VGND VPWR VPWR dadda_fa_4_33_0/B
+ dadda_fa_4_32_1/CIN sky130_fd_sc_hd__fa_2
XU$$3947 U$$3947/A _673_/Q VGND VGND VPWR VPWR U$$3947/X sky130_fd_sc_hd__xor2_1
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$280 final_adder.U$$280/A final_adder.U$$280/B VGND VGND VPWR VPWR
+ final_adder.U$$332/B sky130_fd_sc_hd__and2_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3958 U$$4506/A1 U$$3970/A2 U$$4508/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3959/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$291 final_adder.U$$290/A final_adder.U$$197/X final_adder.U$$199/X
+ VGND VGND VPWR VPWR final_adder.U$$291/X sky130_fd_sc_hd__a21o_1
X_606_ _611_/CLK _606_/D VGND VGND VPWR VPWR _606_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3969 U$$3969/A U$$3969/B VGND VGND VPWR VPWR U$$3969/X sky130_fd_sc_hd__xor2_1
XU$$130 U$$952/A1 U$$4/X U$$952/B1 U$$5/X VGND VGND VPWR VPWR U$$131/A sky130_fd_sc_hd__a22o_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$141 U$$139/Y _618_/Q U$$89/B U$$140/X U$$137/Y VGND VGND VPWR VPWR U$$141/X sky130_fd_sc_hd__a32o_4
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$152 U$$152/A U$$242/B VGND VGND VPWR VPWR U$$152/X sky130_fd_sc_hd__xor2_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$163 _561_/Q U$$141/X U$$987/A1 U$$142/X VGND VGND VPWR VPWR U$$164/A sky130_fd_sc_hd__a22o_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$174 U$$174/A U$$262/B VGND VGND VPWR VPWR U$$174/X sky130_fd_sc_hd__xor2_1
XFILLER_33_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_537_ _537_/CLK _537_/D VGND VGND VPWR VPWR _537_/Q sky130_fd_sc_hd__dfxtp_1
XU$$185 _572_/Q U$$141/X U$$735/A1 U$$142/X VGND VGND VPWR VPWR U$$186/A sky130_fd_sc_hd__a22o_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$196 U$$196/A U$$274/A VGND VGND VPWR VPWR U$$196/X sky130_fd_sc_hd__xor2_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_468_ _480_/CLK _468_/D VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_399_ _543_/CLK _399_/D VGND VGND VPWR VPWR _399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_91_4 dadda_fa_2_91_4/A dadda_fa_2_91_4/B dadda_fa_2_91_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_1/CIN dadda_fa_3_91_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_84_3 dadda_fa_2_84_3/A dadda_fa_2_84_3/B dadda_fa_2_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/B dadda_fa_3_84_3/B sky130_fd_sc_hd__fa_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_77_2 dadda_fa_2_77_2/A dadda_fa_2_77_2/B dadda_fa_2_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/A dadda_fa_3_77_3/A sky130_fd_sc_hd__fa_2
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk _632_/CLK VGND VGND VPWR VPWR _339_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_5_54_1 dadda_fa_5_54_1/A dadda_fa_5_54_1/B dadda_fa_5_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/B dadda_fa_7_54_0/A sky130_fd_sc_hd__fa_2
XFILLER_68_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_47_0 dadda_fa_5_47_0/A dadda_fa_5_47_0/B dadda_fa_5_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/A dadda_fa_6_47_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_100_1 U$$2867/X U$$3000/X U$$3133/X VGND VGND VPWR VPWR dadda_fa_3_101_1/CIN
+ dadda_fa_3_100_3/A sky130_fd_sc_hd__fa_1
XFILLER_36_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_121_0 U$$4372/X U$$4505/X input153/X VGND VGND VPWR VPWR dadda_fa_6_122_0/A
+ dadda_fa_6_121_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_72_1 U$$2412/X U$$2545/X U$$2678/X VGND VGND VPWR VPWR dadda_fa_2_73_0/CIN
+ dadda_fa_2_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_0 U$$2531/X U$$2664/X U$$2797/X VGND VGND VPWR VPWR dadda_fa_2_66_0/B
+ dadda_fa_2_65_3/B sky130_fd_sc_hd__fa_1
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2509 U$$2509/A U$$2533/B VGND VGND VPWR VPWR U$$2509/X sky130_fd_sc_hd__xor2_1
XFILLER_27_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1808 U$$1808/A U$$1856/B VGND VGND VPWR VPWR U$$1808/X sky130_fd_sc_hd__xor2_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1819 _567_/Q U$$1897/A2 U$$3191/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1820/A sky130_fd_sc_hd__a22o_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _448_/CLK _322_/D VGND VGND VPWR VPWR _322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_253_ _503_/CLK _253_/D VGND VGND VPWR VPWR _253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_184_ _329_/CLK _184_/D VGND VGND VPWR VPWR _184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_736__788 VGND VGND VPWR VPWR _736__788/HI U$$2609/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_3_94_2 dadda_fa_3_94_2/A dadda_fa_3_94_2/B dadda_fa_3_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/A dadda_fa_4_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_87_1 dadda_fa_3_87_1/A dadda_fa_3_87_1/B dadda_fa_3_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/CIN dadda_fa_4_87_2/A sky130_fd_sc_hd__fa_2
XFILLER_159_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_64_0 dadda_fa_6_64_0/A dadda_fa_6_64_0/B dadda_fa_6_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_65_0/B dadda_fa_7_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater708 U$$4438/A1 VGND VGND VPWR VPWR U$$54/A1 sky130_fd_sc_hd__buf_12
XFILLER_42_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater719 _571_/Q VGND VGND VPWR VPWR U$$46/A1 sky130_fd_sc_hd__buf_12
XU$$4401 U$$4401/A U$$4401/B VGND VGND VPWR VPWR U$$4401/X sky130_fd_sc_hd__xor2_2
XFILLER_38_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4412 _562_/Q U$$4388/X _563_/Q U$$4389/X VGND VGND VPWR VPWR U$$4413/A sky130_fd_sc_hd__a22o_1
XU$$4423 U$$4423/A U$$4423/B VGND VGND VPWR VPWR U$$4423/X sky130_fd_sc_hd__xor2_4
XFILLER_38_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4434 U$$735/A1 U$$4388/X _574_/Q U$$4389/X VGND VGND VPWR VPWR U$$4435/A sky130_fd_sc_hd__a22o_2
XU$$3700 _670_/Q VGND VGND VPWR VPWR U$$3702/B sky130_fd_sc_hd__inv_1
XU$$4445 U$$4445/A U$$4445/B VGND VGND VPWR VPWR U$$4445/X sky130_fd_sc_hd__xor2_1
XFILLER_49_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4456 U$$70/B1 U$$4388/X U$$759/A1 U$$4389/X VGND VGND VPWR VPWR U$$4457/A sky130_fd_sc_hd__a22o_1
XU$$3711 U$$12/A1 U$$3783/A2 _555_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3712/A sky130_fd_sc_hd__a22o_1
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4467 U$$4467/A U$$4467/B VGND VGND VPWR VPWR U$$4467/X sky130_fd_sc_hd__xor2_4
Xdadda_fa_4_116_1 U$$4229/X U$$4362/X U$$4495/X VGND VGND VPWR VPWR dadda_fa_5_117_0/B
+ dadda_fa_5_116_1/B sky130_fd_sc_hd__fa_2
XU$$3722 U$$3722/A U$$3756/B VGND VGND VPWR VPWR U$$3722/X sky130_fd_sc_hd__xor2_1
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4478 U$$94/A1 U$$4388/X U$$94/B1 U$$4389/X VGND VGND VPWR VPWR U$$4479/A sky130_fd_sc_hd__a22o_1
XU$$3733 _565_/Q U$$3783/A2 U$$4283/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3734/A sky130_fd_sc_hd__a22o_1
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3744 U$$3744/A U$$3794/B VGND VGND VPWR VPWR U$$3744/X sky130_fd_sc_hd__xor2_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4489 U$$4489/A U$$4489/B VGND VGND VPWR VPWR U$$4489/X sky130_fd_sc_hd__xor2_2
Xdadda_fa_4_109_0 dadda_fa_4_109_0/A dadda_fa_4_109_0/B dadda_fa_4_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/A dadda_fa_5_109_1/A sky130_fd_sc_hd__fa_2
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3755 U$$4303/A1 U$$3783/A2 U$$4442/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3756/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3766 U$$3766/A U$$3784/B VGND VGND VPWR VPWR U$$3766/X sky130_fd_sc_hd__xor2_1
XFILLER_80_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3777 _587_/Q U$$3795/A2 U$$765/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3778/A sky130_fd_sc_hd__a22o_1
XFILLER_92_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3788 U$$3788/A _671_/Q VGND VGND VPWR VPWR U$$3788/X sky130_fd_sc_hd__xor2_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3799 U$$4484/A1 U$$3703/X U$$4486/A1 U$$3704/X VGND VGND VPWR VPWR U$$3800/A sky130_fd_sc_hd__a22o_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_82_0 U$$4294/X U$$4427/X input237/X VGND VGND VPWR VPWR dadda_fa_3_83_0/B
+ dadda_fa_3_82_2/B sky130_fd_sc_hd__fa_2
XFILLER_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_685__905 VGND VGND VPWR VPWR _685__905/HI _685__905/LO sky130_fd_sc_hd__conb_1
XFILLER_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_51_6 U$$2503/X U$$2636/X U$$2769/X VGND VGND VPWR VPWR dadda_fa_2_52_2/B
+ dadda_fa_2_51_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_3_0 input190/X dadda_fa_7_3_0/B dadda_ha_6_3_0/SUM VGND VGND VPWR VPWR
+ _428_/D _299_/D sky130_fd_sc_hd__fa_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_81_0 dadda_fa_7_81_0/A dadda_fa_7_81_0/B dadda_fa_7_81_0/CIN VGND VGND
+ VPWR VPWR _506_/D _377_/D sky130_fd_sc_hd__fa_1
XFILLER_109_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_97_0 dadda_fa_4_97_0/A dadda_fa_4_97_0/B dadda_fa_4_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/A dadda_fa_5_97_1/A sky130_fd_sc_hd__fa_1
XFILLER_153_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3007 U$$4514/A1 U$$3009/A2 U$$4379/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$3008/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3018 U$$3016/Y _660_/Q _659_/Q U$$3017/X U$$3014/Y VGND VGND VPWR VPWR U$$3018/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3029 U$$3029/A U$$3085/B VGND VGND VPWR VPWR U$$3029/X sky130_fd_sc_hd__xor2_1
XFILLER_90_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2306 U$$799/A1 U$$2316/A2 U$$938/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2307/A sky130_fd_sc_hd__a22o_1
XU$$2317 U$$2317/A _649_/Q VGND VGND VPWR VPWR U$$2317/X sky130_fd_sc_hd__xor2_1
XFILLER_75_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2328 _649_/Q VGND VGND VPWR VPWR U$$2328/Y sky130_fd_sc_hd__inv_1
XFILLER_90_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2339 _553_/Q U$$2421/A2 U$$4122/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2340/A sky130_fd_sc_hd__a22o_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1605 U$$96/B1 U$$1605/A2 U$$785/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1606/A sky130_fd_sc_hd__a22o_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1616 U$$1616/A U$$1643/A VGND VGND VPWR VPWR U$$1616/X sky130_fd_sc_hd__xor2_1
XU$$1627 U$$4504/A1 U$$1641/A2 U$$944/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1628/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1638 U$$1638/A U$$1643/A VGND VGND VPWR VPWR U$$1638/X sky130_fd_sc_hd__xor2_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1649 U$$1647/B _639_/Q _640_/Q U$$1644/Y VGND VGND VPWR VPWR U$$1649/X sky130_fd_sc_hd__a22o_4
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _331_/CLK _305_/D VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_236_ _499_/CLK _236_/D VGND VGND VPWR VPWR _236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_61_5 dadda_fa_2_61_5/A dadda_fa_2_61_5/B dadda_fa_2_61_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_2/A dadda_fa_4_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_111_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater505 U$$1649/X VGND VGND VPWR VPWR U$$1770/B2 sky130_fd_sc_hd__buf_12
Xrepeater516 _679_/Q VGND VGND VPWR VPWR U$$4332/B sky130_fd_sc_hd__buf_12
Xrepeater527 U$$3794/B VGND VGND VPWR VPWR U$$3784/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_54_4 dadda_fa_2_54_4/A dadda_fa_2_54_4/B dadda_fa_2_54_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/CIN dadda_fa_3_54_3/CIN sky130_fd_sc_hd__fa_2
Xrepeater538 _665_/Q VGND VGND VPWR VPWR U$$3403/B sky130_fd_sc_hd__buf_12
XFILLER_133_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4220 U$$4494/A1 U$$4244/A2 U$$4496/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4221/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4231 U$$4231/A U$$4246/A VGND VGND VPWR VPWR U$$4231/X sky130_fd_sc_hd__xor2_1
XFILLER_65_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater549 U$$2871/B VGND VGND VPWR VPWR U$$2839/B sky130_fd_sc_hd__buf_12
XU$$4242 U$$4379/A1 U$$4244/A2 U$$819/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4243/A
+ sky130_fd_sc_hd__a22o_1
XU$$4253 U$$4253/A1 U$$4251/X U$$4255/A1 U$$4252/X VGND VGND VPWR VPWR U$$4254/A sky130_fd_sc_hd__a22o_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_47_3 dadda_fa_2_47_3/A dadda_fa_2_47_3/B dadda_fa_2_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/B dadda_fa_3_47_3/B sky130_fd_sc_hd__fa_2
XU$$4264 U$$4264/A _679_/Q VGND VGND VPWR VPWR U$$4264/X sky130_fd_sc_hd__xor2_1
XU$$4275 _562_/Q U$$4377/A2 _563_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4276/A sky130_fd_sc_hd__a22o_1
XU$$3530 U$$3530/A U$$3536/B VGND VGND VPWR VPWR U$$3530/X sky130_fd_sc_hd__xor2_1
XU$$4286 U$$4286/A U$$4332/B VGND VGND VPWR VPWR U$$4286/X sky130_fd_sc_hd__xor2_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3541 U$$4500/A1 U$$3429/X U$$4502/A1 U$$3430/X VGND VGND VPWR VPWR U$$3542/A sky130_fd_sc_hd__a22o_1
XU$$3552 U$$3552/A U$$3561/A VGND VGND VPWR VPWR U$$3552/X sky130_fd_sc_hd__xor2_1
XU$$4297 U$$735/A1 U$$4251/X _574_/Q U$$4252/X VGND VGND VPWR VPWR U$$4298/A sky130_fd_sc_hd__a22o_1
XU$$3563 _668_/Q VGND VGND VPWR VPWR U$$3565/B sky130_fd_sc_hd__inv_1
XFILLER_81_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3574 U$$12/A1 U$$3678/A2 _555_/Q U$$3678/B2 VGND VGND VPWR VPWR U$$3575/A sky130_fd_sc_hd__a22o_1
XFILLER_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_17_1 dadda_fa_5_17_1/A dadda_fa_5_17_1/B dadda_fa_5_17_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/B dadda_fa_7_17_0/A sky130_fd_sc_hd__fa_2
XU$$2840 U$$98/B1 U$$2744/X U$$4486/A1 U$$2745/X VGND VGND VPWR VPWR U$$2841/A sky130_fd_sc_hd__a22o_1
XU$$3585 U$$3585/A U$$3625/B VGND VGND VPWR VPWR U$$3585/X sky130_fd_sc_hd__xor2_1
XU$$2851 U$$2851/A U$$2871/B VGND VGND VPWR VPWR U$$2851/X sky130_fd_sc_hd__xor2_1
XU$$3596 _565_/Q U$$3624/A2 _566_/Q U$$3624/B2 VGND VGND VPWR VPWR U$$3597/A sky130_fd_sc_hd__a22o_1
XU$$2862 U$$4506/A1 U$$2744/X U$$4508/A1 U$$2870/B2 VGND VGND VPWR VPWR U$$2863/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2873 U$$2873/A _657_/Q VGND VGND VPWR VPWR U$$2873/X sky130_fd_sc_hd__xor2_1
XU$$2884 U$$2884/A U$$2996/B VGND VGND VPWR VPWR U$$2884/X sky130_fd_sc_hd__xor2_1
XFILLER_179_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2895 U$$4265/A1 U$$3009/A2 U$$979/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2896/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_4_120_1 U$$4237/X U$$4370/X VGND VGND VPWR VPWR dadda_fa_5_121_1/B dadda_ha_4_120_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_43_4 U$$1689/X U$$1822/X VGND VGND VPWR VPWR dadda_fa_2_44_4/A dadda_fa_3_43_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_4_13_2 U$$831/X input161/X VGND VGND VPWR VPWR dadda_fa_5_14_0/CIN dadda_ha_4_13_2/SUM
+ sky130_fd_sc_hd__ha_1
XU$$707 U$$22/A1 U$$689/X _560_/Q U$$817/B2 VGND VGND VPWR VPWR U$$708/A sky130_fd_sc_hd__a22o_1
XFILLER_57_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$718 U$$718/A U$$784/B VGND VGND VPWR VPWR U$$718/X sky130_fd_sc_hd__xor2_1
XFILLER_72_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$729 _570_/Q U$$689/X U$$46/A1 U$$817/B2 VGND VGND VPWR VPWR U$$730/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_2 U$$889/X U$$1022/X U$$1155/X VGND VGND VPWR VPWR dadda_fa_2_43_3/CIN
+ dadda_fa_2_42_5/B sky130_fd_sc_hd__fa_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_12_0 U$$31/X U$$164/X U$$297/X VGND VGND VPWR VPWR dadda_fa_5_13_0/A dadda_fa_5_12_1/A
+ sky130_fd_sc_hd__fa_2
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_64_3 dadda_fa_3_64_3/A dadda_fa_3_64_3/B dadda_fa_3_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/B dadda_fa_4_64_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_57_2 dadda_fa_3_57_2/A dadda_fa_3_57_2/B dadda_fa_3_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/A dadda_fa_4_57_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_27_0 dadda_fa_6_27_0/A dadda_fa_6_27_0/B dadda_fa_6_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_28_0/B dadda_fa_7_27_0/CIN sky130_fd_sc_hd__fa_1
XU$$2103 U$$48/A1 U$$2117/A2 U$$50/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2104/A sky130_fd_sc_hd__a22o_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2114 U$$2114/A U$$2118/B VGND VGND VPWR VPWR U$$2114/X sky130_fd_sc_hd__xor2_1
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2125 U$$68/B1 U$$2161/A2 U$$72/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2126/A sky130_fd_sc_hd__a22o_1
XU$$2136 U$$2136/A U$$2186/B VGND VGND VPWR VPWR U$$2136/X sky130_fd_sc_hd__xor2_1
XU$$2147 _594_/Q U$$2189/A2 _595_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2148/A sky130_fd_sc_hd__a22o_1
XFILLER_62_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1402 U$$30/B1 U$$1474/A2 U$$3457/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1403/A sky130_fd_sc_hd__a22o_1
XU$$2158 U$$2158/A U$$2192/A VGND VGND VPWR VPWR U$$2158/X sky130_fd_sc_hd__xor2_1
XU$$1413 U$$1413/A U$$1461/B VGND VGND VPWR VPWR U$$1413/X sky130_fd_sc_hd__xor2_1
XU$$1424 U$$876/A1 U$$1472/A2 U$$878/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1425/A sky130_fd_sc_hd__a22o_1
XFILLER_90_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2169 U$$799/A1 U$$2189/A2 _606_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2170/A sky130_fd_sc_hd__a22o_1
XU$$1435 U$$1435/A U$$1461/B VGND VGND VPWR VPWR U$$1435/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1446 U$$2953/A1 U$$1472/A2 U$$76/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1447/A sky130_fd_sc_hd__a22o_1
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1457 U$$1457/A U$$1461/B VGND VGND VPWR VPWR U$$1457/X sky130_fd_sc_hd__xor2_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1468 U$$98/A1 U$$1474/A2 U$$98/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1469/A sky130_fd_sc_hd__a22o_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1479 U$$1479/A U$$1479/B VGND VGND VPWR VPWR U$$1479/X sky130_fd_sc_hd__xor2_1
XFILLER_96_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_219_ _474_/CLK _219_/D VGND VGND VPWR VPWR _219_/Q sky130_fd_sc_hd__dfxtp_1
X_751__803 VGND VGND VPWR VPWR _751__803/HI U$$3559/B1 sky130_fd_sc_hd__conb_1
XFILLER_117_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_1_clk clkbuf_1_1_1_clk/A VGND VGND VPWR VPWR clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
Xfinal_adder.U$$109 _533_/Q _405_/Q VGND VGND VPWR VPWR final_adder.U$$237/B1 final_adder.U$$731/A
+ sky130_fd_sc_hd__ha_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_52_1 dadda_fa_2_52_1/A dadda_fa_2_52_1/B dadda_fa_2_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/CIN dadda_fa_3_52_2/CIN sky130_fd_sc_hd__fa_1
XU$$4050 U$$4050/A U$$4109/A VGND VGND VPWR VPWR U$$4050/X sky130_fd_sc_hd__xor2_1
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_45_0 U$$2358/X U$$2491/X U$$2624/X VGND VGND VPWR VPWR dadda_fa_3_46_0/B
+ dadda_fa_3_45_2/B sky130_fd_sc_hd__fa_2
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4061 U$$771/B1 U$$4107/A2 _593_/Q U$$4107/B2 VGND VGND VPWR VPWR U$$4062/A sky130_fd_sc_hd__a22o_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4072 U$$4072/A U$$4109/A VGND VGND VPWR VPWR U$$4072/X sky130_fd_sc_hd__xor2_1
XFILLER_26_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4083 U$$4494/A1 U$$4107/A2 U$$4496/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4084/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4094 U$$4094/A U$$4109/A VGND VGND VPWR VPWR U$$4094/X sky130_fd_sc_hd__xor2_1
XU$$3360 U$$892/B1 U$$3396/A2 U$$4045/B1 U$$3396/B2 VGND VGND VPWR VPWR U$$3361/A
+ sky130_fd_sc_hd__a22o_1
XU$$3371 U$$3371/A U$$3413/B VGND VGND VPWR VPWR U$$3371/X sky130_fd_sc_hd__xor2_1
XU$$3382 _595_/Q U$$3292/X _596_/Q U$$3293/X VGND VGND VPWR VPWR U$$3383/A sky130_fd_sc_hd__a22o_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3393 U$$3393/A U$$3397/B VGND VGND VPWR VPWR U$$3393/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2670 U$$2670/A U$$2694/B VGND VGND VPWR VPWR U$$2670/X sky130_fd_sc_hd__xor2_1
XU$$2681 _587_/Q U$$2607/X _588_/Q U$$2608/X VGND VGND VPWR VPWR U$$2682/A sky130_fd_sc_hd__a22o_1
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2692 U$$2692/A U$$2710/B VGND VGND VPWR VPWR U$$2692/X sky130_fd_sc_hd__xor2_1
XFILLER_34_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1980 U$$4446/A1 U$$2048/A2 U$$3900/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1981/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1991 U$$1991/A U$$1991/B VGND VGND VPWR VPWR U$$1991/X sky130_fd_sc_hd__xor2_1
XFILLER_193_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_74_2 dadda_fa_4_74_2/A dadda_fa_4_74_2/B dadda_fa_4_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/CIN dadda_fa_5_74_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_67_1 dadda_fa_4_67_1/A dadda_fa_4_67_1/B dadda_fa_4_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/B dadda_fa_5_67_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput105 b[46] VGND VGND VPWR VPWR _598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput116 b[56] VGND VGND VPWR VPWR _608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_44_0 dadda_fa_7_44_0/A dadda_fa_7_44_0/B dadda_fa_7_44_0/CIN VGND VGND
+ VPWR VPWR _469_/D _340_/D sky130_fd_sc_hd__fa_2
XFILLER_131_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput127 b[8] VGND VGND VPWR VPWR _560_/D sky130_fd_sc_hd__clkbuf_4
Xinput138 c[108] VGND VGND VPWR VPWR input138/X sky130_fd_sc_hd__clkbuf_2
Xdadda_ha_1_34_0 U$$75/X U$$208/X VGND VGND VPWR VPWR dadda_fa_2_35_5/CIN dadda_fa_3_34_0/A
+ sky130_fd_sc_hd__ha_1
Xinput149 c[118] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$621 final_adder.U$$748/A final_adder.U$$748/B final_adder.U$$621/B1
+ VGND VGND VPWR VPWR final_adder.U$$749/B sky130_fd_sc_hd__a21o_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$632 final_adder.U$$632/A final_adder.U$$632/B VGND VGND VPWR VPWR
+ _178_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$643 final_adder.U$$643/A final_adder.U$$643/B VGND VGND VPWR VPWR
+ _189_/D sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$654 final_adder.U$$654/A final_adder.U$$654/B VGND VGND VPWR VPWR
+ _200_/D sky130_fd_sc_hd__xor2_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$665 final_adder.U$$665/A final_adder.U$$665/B VGND VGND VPWR VPWR
+ _211_/D sky130_fd_sc_hd__xor2_1
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$504 U$$504/A U$$547/A VGND VGND VPWR VPWR U$$504/X sky130_fd_sc_hd__xor2_1
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$676 final_adder.U$$676/A final_adder.U$$676/B VGND VGND VPWR VPWR
+ _222_/D sky130_fd_sc_hd__xor2_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$515 U$$926/A1 U$$545/A2 U$$928/A1 U$$416/X VGND VGND VPWR VPWR U$$516/A sky130_fd_sc_hd__a22o_1
X_570_ _576_/CLK _570_/D VGND VGND VPWR VPWR _570_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$687 final_adder.U$$687/A final_adder.U$$687/B VGND VGND VPWR VPWR
+ _233_/D sky130_fd_sc_hd__xor2_1
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$526 U$$526/A U$$547/A VGND VGND VPWR VPWR U$$526/X sky130_fd_sc_hd__xor2_1
XFILLER_99_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$698 final_adder.U$$698/A final_adder.U$$698/B VGND VGND VPWR VPWR
+ _244_/D sky130_fd_sc_hd__xor2_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$537 U$$948/A1 U$$415/X U$$539/A1 U$$416/X VGND VGND VPWR VPWR U$$538/A sky130_fd_sc_hd__a22o_1
XFILLER_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$548 _623_/Q VGND VGND VPWR VPWR U$$548/Y sky130_fd_sc_hd__inv_1
XFILLER_56_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$559 U$$559/A U$$623/B VGND VGND VPWR VPWR U$$559/X sky130_fd_sc_hd__xor2_1
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_62_0 dadda_fa_3_62_0/A dadda_fa_3_62_0/B dadda_fa_3_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/B dadda_fa_4_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_9_0 U$$25/X U$$158/X VGND VGND VPWR VPWR dadda_fa_5_10_1/A dadda_ha_4_9_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1210 U$$799/A1 U$$1100/X U$$938/A1 U$$1101/X VGND VGND VPWR VPWR U$$1211/A sky130_fd_sc_hd__a22o_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1221 U$$1221/A U$$1232/A VGND VGND VPWR VPWR U$$1221/X sky130_fd_sc_hd__xor2_1
XFILLER_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1232 U$$1232/A VGND VGND VPWR VPWR U$$1232/Y sky130_fd_sc_hd__inv_1
XFILLER_189_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1243 U$$8/B1 U$$1237/X U$$971/A1 U$$1238/X VGND VGND VPWR VPWR U$$1244/A sky130_fd_sc_hd__a22o_1
XFILLER_50_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1254 U$$1254/A U$$1336/B VGND VGND VPWR VPWR U$$1254/X sky130_fd_sc_hd__xor2_1
XU$$1265 U$$32/A1 U$$1237/X U$$34/A1 U$$1238/X VGND VGND VPWR VPWR U$$1266/A sky130_fd_sc_hd__a22o_1
XU$$1276 U$$1276/A U$$1342/B VGND VGND VPWR VPWR U$$1276/X sky130_fd_sc_hd__xor2_1
XU$$1287 U$$54/A1 U$$1237/X U$$56/A1 U$$1238/X VGND VGND VPWR VPWR U$$1288/A sky130_fd_sc_hd__a22o_1
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1298 U$$1298/A U$$1342/B VGND VGND VPWR VPWR U$$1298/X sky130_fd_sc_hd__xor2_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_175_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_84_1 dadda_fa_5_84_1/A dadda_fa_5_84_1/B dadda_fa_5_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/B dadda_fa_7_84_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_77_0 dadda_fa_5_77_0/A dadda_fa_5_77_0/B dadda_fa_5_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/A dadda_fa_6_77_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_76_8 dadda_fa_1_76_8/A dadda_fa_1_76_8/B dadda_fa_1_76_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_77_3/A dadda_fa_3_76_0/A sky130_fd_sc_hd__fa_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_7 dadda_fa_1_69_7/A dadda_fa_1_69_7/B dadda_fa_1_69_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/CIN dadda_fa_2_69_5/CIN sky130_fd_sc_hd__fa_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3190 U$$3190/A U$$3224/B VGND VGND VPWR VPWR U$$3190/X sky130_fd_sc_hd__xor2_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_95_0 U$$2191/Y U$$2325/X U$$2458/X VGND VGND VPWR VPWR dadda_fa_2_96_5/CIN
+ dadda_fa_3_95_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_3_100_3 dadda_fa_3_100_3/A dadda_fa_3_100_3/B dadda_fa_3_100_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/B dadda_fa_4_100_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_2_108_0 _706__926/HI U$$3149/X VGND VGND VPWR VPWR dadda_fa_4_109_0/A dadda_fa_4_108_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_190_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$451 final_adder.U$$274/B final_adder.U$$658/B final_adder.U$$165/X
+ VGND VGND VPWR VPWR final_adder.U$$660/B sky130_fd_sc_hd__a21o_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ _622_/CLK _622_/D VGND VGND VPWR VPWR _622_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$301 U$$301/A U$$357/B VGND VGND VPWR VPWR U$$301/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_107_0 dadda_fa_6_107_0/A dadda_fa_6_107_0/B dadda_fa_6_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_108_0/B dadda_fa_7_107_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_85_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$473 final_adder.U$$296/B final_adder.U$$702/B final_adder.U$$209/X
+ VGND VGND VPWR VPWR final_adder.U$$704/B sky130_fd_sc_hd__a21o_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$312 U$$38/A1 U$$278/X U$$40/A1 U$$279/X VGND VGND VPWR VPWR U$$313/A sky130_fd_sc_hd__a22o_1
XFILLER_85_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$323 U$$323/A U$$391/B VGND VGND VPWR VPWR U$$323/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$495 final_adder.U$$252/X final_adder.U$$746/B final_adder.U$$253/X
+ VGND VGND VPWR VPWR final_adder.U$$748/B sky130_fd_sc_hd__a21o_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$334 U$$60/A1 U$$278/X U$$62/A1 U$$279/X VGND VGND VPWR VPWR U$$335/A sky130_fd_sc_hd__a22o_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$345 U$$345/A U$$357/B VGND VGND VPWR VPWR U$$345/X sky130_fd_sc_hd__xor2_1
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_553_ _573_/CLK _553_/D VGND VGND VPWR VPWR _553_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$356 U$$82/A1 U$$278/X U$$84/A1 U$$279/X VGND VGND VPWR VPWR U$$357/A sky130_fd_sc_hd__a22o_1
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$367 U$$367/A _621_/Q VGND VGND VPWR VPWR U$$367/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_27_3 dadda_fa_3_27_3/A dadda_fa_3_27_3/B dadda_fa_3_27_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_28_1/B dadda_fa_4_27_2/CIN sky130_fd_sc_hd__fa_2
XU$$378 U$$926/A1 U$$278/X U$$928/A1 U$$279/X VGND VGND VPWR VPWR U$$379/A sky130_fd_sc_hd__a22o_1
XFILLER_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$389 U$$389/A _621_/Q VGND VGND VPWR VPWR U$$389/X sky130_fd_sc_hd__xor2_1
XFILLER_83_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_484_ _499_/CLK _484_/D VGND VGND VPWR VPWR _484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_94_0 dadda_fa_6_94_0/A dadda_fa_6_94_0/B dadda_fa_6_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_95_0/B dadda_fa_7_94_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$890 U$$68/A1 U$$910/A2 U$$68/B1 U$$910/B2 VGND VGND VPWR VPWR U$$891/A sky130_fd_sc_hd__a22o_1
XU$$1040 U$$1040/A U$$980/B VGND VGND VPWR VPWR U$$1040/X sky130_fd_sc_hd__xor2_1
XU$$1051 U$$914/A1 U$$1093/A2 U$$92/B1 U$$1073/B2 VGND VGND VPWR VPWR U$$1052/A sky130_fd_sc_hd__a22o_1
XU$$1062 U$$1062/A U$$980/B VGND VGND VPWR VPWR U$$1062/X sky130_fd_sc_hd__xor2_1
XU$$1073 U$$799/A1 U$$1093/A2 U$$938/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1074/A sky130_fd_sc_hd__a22o_1
XU$$1084 U$$1084/A _631_/Q VGND VGND VPWR VPWR U$$1084/X sky130_fd_sc_hd__xor2_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1095 _631_/Q VGND VGND VPWR VPWR U$$1095/Y sky130_fd_sc_hd__inv_1
XFILLER_137_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_81_6 U$$3627/X U$$3760/X U$$3893/X VGND VGND VPWR VPWR dadda_fa_2_82_3/A
+ dadda_fa_2_81_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_74_5 U$$3746/X U$$3879/X U$$4012/X VGND VGND VPWR VPWR dadda_fa_2_75_2/A
+ dadda_fa_2_74_5/A sky130_fd_sc_hd__fa_2
XFILLER_113_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_4 U$$4131/X U$$4264/X U$$4397/X VGND VGND VPWR VPWR dadda_fa_2_68_1/CIN
+ dadda_fa_2_67_4/CIN sky130_fd_sc_hd__fa_2
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_37_2 dadda_fa_4_37_2/A dadda_fa_4_37_2/B dadda_fa_4_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/CIN dadda_fa_5_37_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_63_5 U$$2128/X U$$2261/X VGND VGND VPWR VPWR dadda_fa_1_64_7/A dadda_fa_2_63_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_162_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_3 U$$1328/X U$$1461/X U$$1594/X VGND VGND VPWR VPWR dadda_fa_1_63_6/B
+ dadda_fa_1_62_8/B sky130_fd_sc_hd__fa_1
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3904 U$$4178/A1 U$$3912/A2 U$$70/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3905/A sky130_fd_sc_hd__a22o_1
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3915 U$$3915/A U$$3969/B VGND VGND VPWR VPWR U$$3915/X sky130_fd_sc_hd__xor2_1
XFILLER_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3926 _593_/Q U$$3970/A2 U$$4476/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3927/A sky130_fd_sc_hd__a22o_1
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3937 U$$3937/A _673_/Q VGND VGND VPWR VPWR U$$3937/X sky130_fd_sc_hd__xor2_1
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$270 final_adder.U$$270/A final_adder.U$$270/B VGND VGND VPWR VPWR
+ final_adder.U$$326/A sky130_fd_sc_hd__and2_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3948 U$$4496/A1 U$$3970/A2 U$$936/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3949/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$281 final_adder.U$$280/A final_adder.U$$177/X final_adder.U$$179/X
+ VGND VGND VPWR VPWR final_adder.U$$281/X sky130_fd_sc_hd__a21o_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_32_1 dadda_fa_3_32_1/A dadda_fa_3_32_1/B dadda_fa_3_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_0/CIN dadda_fa_4_32_2/A sky130_fd_sc_hd__fa_2
XU$$120 _608_/Q U$$4/X _609_/Q U$$5/X VGND VGND VPWR VPWR U$$121/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$292 final_adder.U$$292/A final_adder.U$$292/B VGND VGND VPWR VPWR
+ final_adder.U$$338/B sky130_fd_sc_hd__and2_1
X_605_ _611_/CLK _605_/D VGND VGND VPWR VPWR _605_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3959 U$$3959/A _673_/Q VGND VGND VPWR VPWR U$$3959/X sky130_fd_sc_hd__xor2_1
XU$$131 U$$131/A _617_/Q VGND VGND VPWR VPWR U$$131/X sky130_fd_sc_hd__xor2_1
XFILLER_40_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$142 U$$140/B U$$89/B _618_/Q U$$137/Y VGND VGND VPWR VPWR U$$142/X sky130_fd_sc_hd__a22o_4
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$153 U$$16/A1 U$$141/X U$$18/A1 U$$142/X VGND VGND VPWR VPWR U$$154/A sky130_fd_sc_hd__a22o_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_25_0 U$$722/X U$$855/X U$$988/X VGND VGND VPWR VPWR dadda_fa_4_26_0/B
+ dadda_fa_4_25_1/CIN sky130_fd_sc_hd__fa_1
XU$$164 U$$164/A U$$242/B VGND VGND VPWR VPWR U$$164/X sky130_fd_sc_hd__xor2_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$175 U$$38/A1 U$$141/X U$$40/A1 U$$142/X VGND VGND VPWR VPWR U$$176/A sky130_fd_sc_hd__a22o_1
X_536_ _536_/CLK _536_/D VGND VGND VPWR VPWR _536_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$186 U$$186/A U$$262/B VGND VGND VPWR VPWR U$$186/X sky130_fd_sc_hd__xor2_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$197 U$$60/A1 U$$141/X U$$62/A1 U$$142/X VGND VGND VPWR VPWR U$$198/A sky130_fd_sc_hd__a22o_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_467_ _467_/CLK _467_/D VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_398_ _527_/CLK _398_/D VGND VGND VPWR VPWR _398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_91_5 dadda_fa_2_91_5/A dadda_fa_2_91_5/B dadda_fa_2_91_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_2/A dadda_fa_4_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_84_4 dadda_fa_2_84_4/A dadda_fa_2_84_4/B dadda_fa_2_84_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/CIN dadda_fa_3_84_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_77_3 dadda_fa_2_77_3/A dadda_fa_2_77_3/B dadda_fa_2_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/B dadda_fa_3_77_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_47_1 dadda_fa_5_47_1/A dadda_fa_5_47_1/B dadda_fa_5_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/B dadda_fa_7_47_0/A sky130_fd_sc_hd__fa_2
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_100_2 U$$3266/X U$$3399/X U$$3532/X VGND VGND VPWR VPWR dadda_fa_3_101_2/A
+ dadda_fa_3_100_3/B sky130_fd_sc_hd__fa_1
XFILLER_51_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_121_1 dadda_fa_5_121_1/A dadda_fa_5_121_1/B dadda_fa_5_121_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_122_0/B dadda_fa_7_121_0/A sky130_fd_sc_hd__fa_2
XFILLER_20_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_114_0 dadda_fa_5_114_0/A dadda_fa_5_114_0/B dadda_fa_5_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/A dadda_fa_6_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_1_72_2 U$$2811/X U$$2944/X U$$3077/X VGND VGND VPWR VPWR dadda_fa_2_73_1/A
+ dadda_fa_2_72_4/A sky130_fd_sc_hd__fa_2
XFILLER_63_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_1 U$$2930/X U$$3063/X U$$3196/X VGND VGND VPWR VPWR dadda_fa_2_66_0/CIN
+ dadda_fa_2_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_42_0 dadda_fa_4_42_0/A dadda_fa_4_42_0/B dadda_fa_4_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/A dadda_fa_5_42_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_58_0 U$$1586/X U$$1719/X U$$1852/X VGND VGND VPWR VPWR dadda_fa_2_59_0/B
+ dadda_fa_2_58_3/B sky130_fd_sc_hd__fa_2
XFILLER_86_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1809 U$$987/A1 U$$1867/A2 U$$28/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1810/A sky130_fd_sc_hd__a22o_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_321_ _448_/CLK _321_/D VGND VGND VPWR VPWR _321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_252_ _503_/CLK _252_/D VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_183_ _464_/CLK _183_/D VGND VGND VPWR VPWR _183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_94_3 dadda_fa_3_94_3/A dadda_fa_3_94_3/B dadda_fa_3_94_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/B dadda_fa_4_94_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_87_2 dadda_fa_3_87_2/A dadda_fa_3_87_2/B dadda_fa_3_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/A dadda_fa_4_87_2/B sky130_fd_sc_hd__fa_1
XFILLER_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_0_54_1 U$$514/X U$$647/X VGND VGND VPWR VPWR dadda_fa_1_55_8/B dadda_fa_2_54_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_6_57_0 dadda_fa_6_57_0/A dadda_fa_6_57_0/B dadda_fa_6_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_58_0/B dadda_fa_7_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater709 _575_/Q VGND VGND VPWR VPWR U$$4438/A1 sky130_fd_sc_hd__buf_12
XU$$4402 _557_/Q U$$4388/X _558_/Q U$$4389/X VGND VGND VPWR VPWR U$$4403/A sky130_fd_sc_hd__a22o_1
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4413 U$$4413/A U$$4413/B VGND VGND VPWR VPWR U$$4413/X sky130_fd_sc_hd__xor2_2
XU$$4424 U$$4424/A1 U$$4388/X _569_/Q U$$4389/X VGND VGND VPWR VPWR U$$4425/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_60_0 U$$127/X U$$260/X U$$393/X VGND VGND VPWR VPWR dadda_fa_1_61_6/A
+ dadda_fa_1_60_7/CIN sky130_fd_sc_hd__fa_2
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4435 U$$4435/A U$$4435/B VGND VGND VPWR VPWR U$$4435/X sky130_fd_sc_hd__xor2_4
XU$$4446 U$$4446/A1 U$$4388/X _580_/Q U$$4389/X VGND VGND VPWR VPWR U$$4447/A sky130_fd_sc_hd__a22o_1
XFILLER_92_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3701 _671_/Q VGND VGND VPWR VPWR U$$3701/Y sky130_fd_sc_hd__inv_1
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3712 U$$3712/A U$$3784/B VGND VGND VPWR VPWR U$$3712/X sky130_fd_sc_hd__xor2_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_116_2 input147/X dadda_fa_4_116_2/B dadda_ha_3_116_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_5_117_0/CIN dadda_fa_5_116_1/CIN sky130_fd_sc_hd__fa_1
XU$$4457 U$$4457/A U$$4457/B VGND VGND VPWR VPWR U$$4457/X sky130_fd_sc_hd__xor2_1
XFILLER_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4468 U$$632/A1 U$$4388/X U$$771/A1 U$$4389/X VGND VGND VPWR VPWR U$$4469/A sky130_fd_sc_hd__a22o_1
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3723 U$$983/A1 U$$3783/A2 U$$4273/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3724/A
+ sky130_fd_sc_hd__a22o_1
XU$$4479 U$$4479/A U$$4479/B VGND VGND VPWR VPWR U$$4479/X sky130_fd_sc_hd__xor2_2
XU$$3734 U$$3734/A U$$3756/B VGND VGND VPWR VPWR U$$3734/X sky130_fd_sc_hd__xor2_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3745 _571_/Q U$$3783/A2 _572_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3746/A sky130_fd_sc_hd__a22o_1
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3756 U$$3756/A U$$3756/B VGND VGND VPWR VPWR U$$3756/X sky130_fd_sc_hd__xor2_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_109_1 dadda_fa_4_109_1/A dadda_fa_4_109_1/B dadda_fa_4_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/B dadda_fa_5_109_1/B sky130_fd_sc_hd__fa_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3767 _582_/Q U$$3783/A2 U$$70/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3768/A sky130_fd_sc_hd__a22o_1
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3778 U$$3778/A _671_/Q VGND VGND VPWR VPWR U$$3778/X sky130_fd_sc_hd__xor2_1
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3789 _593_/Q U$$3795/A2 _594_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3790/A sky130_fd_sc_hd__a22o_1
XFILLER_79_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_519_ _535_/CLK _519_/D VGND VGND VPWR VPWR _519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_82_1 dadda_fa_2_82_1/A dadda_fa_2_82_1/B dadda_fa_2_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_0/CIN dadda_fa_3_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_75_0 dadda_fa_2_75_0/A dadda_fa_2_75_0/B dadda_fa_2_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/B dadda_fa_3_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_141_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_51_7 U$$2902/X U$$3035/X U$$3168/X VGND VGND VPWR VPWR dadda_fa_2_52_2/CIN
+ dadda_fa_2_51_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_97_1 dadda_fa_4_97_1/A dadda_fa_4_97_1/B dadda_fa_4_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/B dadda_fa_5_97_1/B sky130_fd_sc_hd__fa_1
XFILLER_153_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_74_0 dadda_fa_7_74_0/A dadda_fa_7_74_0/B dadda_fa_7_74_0/CIN VGND VGND
+ VPWR VPWR _499_/D _370_/D sky130_fd_sc_hd__fa_1
XFILLER_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3008 U$$3008/A _659_/Q VGND VGND VPWR VPWR U$$3008/X sky130_fd_sc_hd__xor2_1
XFILLER_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3019 U$$3017/B _659_/Q _660_/Q U$$3014/Y VGND VGND VPWR VPWR U$$3019/X sky130_fd_sc_hd__a22o_4
XFILLER_74_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2307 U$$2307/A U$$2327/B VGND VGND VPWR VPWR U$$2307/X sky130_fd_sc_hd__xor2_1
XU$$2318 U$$4510/A1 U$$2326/A2 _612_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2319/A sky130_fd_sc_hd__a22o_1
XU$$2329 _649_/Q VGND VGND VPWR VPWR U$$2329/Y sky130_fd_sc_hd__inv_1
XFILLER_15_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1606 U$$1606/A U$$1643/A VGND VGND VPWR VPWR U$$1606/X sky130_fd_sc_hd__xor2_1
XU$$1617 _603_/Q U$$1641/A2 _604_/Q U$$1641/B2 VGND VGND VPWR VPWR U$$1618/A sky130_fd_sc_hd__a22o_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1628 U$$1628/A _639_/Q VGND VGND VPWR VPWR U$$1628/X sky130_fd_sc_hd__xor2_1
XFILLER_15_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1639 U$$952/B1 U$$1641/A2 U$$956/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1640/A sky130_fd_sc_hd__a22o_1
XFILLER_72_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _465_/CLK _304_/D VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ _499_/CLK hold1/X VGND VGND VPWR VPWR _235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_92_0 dadda_fa_3_92_0/A dadda_fa_3_92_0/B dadda_fa_3_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/B dadda_fa_4_92_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater506 U$$1591/B2 VGND VGND VPWR VPWR U$$1605/B2 sky130_fd_sc_hd__buf_12
Xrepeater517 _677_/Q VGND VGND VPWR VPWR U$$4246/A sky130_fd_sc_hd__buf_12
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4210 U$$4484/A1 U$$4244/A2 U$$4486/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4211/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater528 U$$3794/B VGND VGND VPWR VPWR U$$3835/A sky130_fd_sc_hd__buf_12
Xdadda_fa_2_54_5 dadda_fa_2_54_5/A dadda_fa_2_54_5/B dadda_fa_2_54_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_2/A dadda_fa_4_54_0/A sky130_fd_sc_hd__fa_1
XU$$4221 U$$4221/A U$$4246/A VGND VGND VPWR VPWR U$$4221/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_121_0 U$$3972/Y U$$4106/X U$$4239/X VGND VGND VPWR VPWR dadda_fa_5_122_1/B
+ dadda_fa_5_121_1/CIN sky130_fd_sc_hd__fa_1
Xrepeater539 _663_/Q VGND VGND VPWR VPWR U$$3224/B sky130_fd_sc_hd__buf_12
XFILLER_120_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4232 U$$4506/A1 U$$4244/A2 U$$4508/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4233/A
+ sky130_fd_sc_hd__a22o_1
XU$$4243 U$$4243/A U$$4246/A VGND VGND VPWR VPWR U$$4243/X sky130_fd_sc_hd__xor2_1
XFILLER_65_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4254 U$$4254/A U$$4332/B VGND VGND VPWR VPWR U$$4254/X sky130_fd_sc_hd__xor2_1
XU$$3520 U$$3520/A U$$3561/A VGND VGND VPWR VPWR U$$3520/X sky130_fd_sc_hd__xor2_1
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_47_4 dadda_fa_2_47_4/A dadda_fa_2_47_4/B dadda_fa_2_47_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/CIN dadda_fa_3_47_3/CIN sky130_fd_sc_hd__fa_2
XU$$4265 U$$4265/A1 U$$4251/X U$$842/A1 U$$4252/X VGND VGND VPWR VPWR U$$4266/A sky130_fd_sc_hd__a22o_1
XU$$4276 U$$4276/A U$$4384/A VGND VGND VPWR VPWR U$$4276/X sky130_fd_sc_hd__xor2_1
XU$$3531 _601_/Q U$$3545/A2 U$$928/B1 U$$3545/B2 VGND VGND VPWR VPWR U$$3532/A sky130_fd_sc_hd__a22o_1
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3542 U$$3542/A U$$3561/A VGND VGND VPWR VPWR U$$3542/X sky130_fd_sc_hd__xor2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4287 U$$4424/A1 U$$4377/A2 _569_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4288/A sky130_fd_sc_hd__a22o_1
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3553 U$$539/A1 U$$3429/X _613_/Q U$$3430/X VGND VGND VPWR VPWR U$$3554/A sky130_fd_sc_hd__a22o_1
XU$$4298 U$$4298/A U$$4332/B VGND VGND VPWR VPWR U$$4298/X sky130_fd_sc_hd__xor2_1
XU$$3564 _669_/Q VGND VGND VPWR VPWR U$$3564/Y sky130_fd_sc_hd__inv_1
XFILLER_34_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3575 U$$3575/A U$$3698/A VGND VGND VPWR VPWR U$$3575/X sky130_fd_sc_hd__xor2_1
XU$$2830 _593_/Q U$$2868/A2 U$$914/A1 U$$2870/B2 VGND VGND VPWR VPWR U$$2831/A sky130_fd_sc_hd__a22o_1
XU$$2841 U$$2841/A _657_/Q VGND VGND VPWR VPWR U$$2841/X sky130_fd_sc_hd__xor2_1
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3586 U$$4271/A1 U$$3624/A2 U$$4273/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3587/A
+ sky130_fd_sc_hd__a22o_1
XU$$2852 U$$934/A1 U$$2868/A2 _605_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2853/A sky130_fd_sc_hd__a22o_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3597 U$$3597/A _669_/Q VGND VGND VPWR VPWR U$$3597/X sky130_fd_sc_hd__xor2_1
XU$$2863 U$$2863/A _657_/Q VGND VGND VPWR VPWR U$$2863/X sky130_fd_sc_hd__xor2_1
XU$$2874 U$$956/A1 U$$2744/X U$$2874/B1 U$$2745/X VGND VGND VPWR VPWR U$$2875/A sky130_fd_sc_hd__a22o_1
XU$$2885 U$$8/A1 U$$3009/A2 U$$8/B1 U$$3009/B2 VGND VGND VPWR VPWR U$$2886/A sky130_fd_sc_hd__a22o_1
XFILLER_179_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2896 U$$2896/A U$$2996/B VGND VGND VPWR VPWR U$$2896/X sky130_fd_sc_hd__xor2_1
XFILLER_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$708 U$$708/A U$$784/B VGND VGND VPWR VPWR U$$708/X sky130_fd_sc_hd__xor2_1
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$719 U$$34/A1 U$$785/A2 U$$36/A1 U$$785/B2 VGND VGND VPWR VPWR U$$720/A sky130_fd_sc_hd__a22o_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_42_3 U$$1288/X U$$1421/X U$$1554/X VGND VGND VPWR VPWR dadda_fa_2_43_4/A
+ dadda_fa_2_42_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_12_1 U$$430/X U$$563/X U$$696/X VGND VGND VPWR VPWR dadda_fa_5_13_0/B
+ dadda_fa_5_12_1/B sky130_fd_sc_hd__fa_1
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_109_0 U$$3150/Y U$$3284/X U$$3417/X VGND VGND VPWR VPWR dadda_fa_4_110_0/B
+ dadda_fa_4_109_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_57_3 dadda_fa_3_57_3/A dadda_fa_3_57_3/B dadda_fa_3_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/B dadda_fa_4_57_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2104 U$$2104/A U$$2118/B VGND VGND VPWR VPWR U$$2104/X sky130_fd_sc_hd__xor2_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2115 U$$4170/A1 U$$2117/A2 U$$3624/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2116/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2126 U$$2126/A _647_/Q VGND VGND VPWR VPWR U$$2126/X sky130_fd_sc_hd__xor2_1
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2137 U$$902/B1 U$$2161/A2 U$$84/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2138/A sky130_fd_sc_hd__a22o_1
XU$$2148 U$$2148/A _647_/Q VGND VGND VPWR VPWR U$$2148/X sky130_fd_sc_hd__xor2_1
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1403 U$$1403/A U$$1461/B VGND VGND VPWR VPWR U$$1403/X sky130_fd_sc_hd__xor2_1
XU$$2159 U$$787/B1 U$$2161/A2 U$$654/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2160/A sky130_fd_sc_hd__a22o_1
XU$$1414 U$$4291/A1 U$$1472/A2 U$$868/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1415/A
+ sky130_fd_sc_hd__a22o_1
XU$$1425 U$$1425/A U$$1505/B VGND VGND VPWR VPWR U$$1425/X sky130_fd_sc_hd__xor2_1
XU$$1436 U$$66/A1 U$$1474/A2 U$$68/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1437/A sky130_fd_sc_hd__a22o_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1447 U$$1447/A U$$1505/B VGND VGND VPWR VPWR U$$1447/X sky130_fd_sc_hd__xor2_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1458 U$$88/A1 U$$1472/A2 U$$90/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1459/A sky130_fd_sc_hd__a22o_1
XFILLER_128_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1469 U$$1469/A U$$1479/B VGND VGND VPWR VPWR U$$1469/X sky130_fd_sc_hd__xor2_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_218_ _480_/CLK _218_/D VGND VGND VPWR VPWR _218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_790__842 VGND VGND VPWR VPWR _790__842/HI U$$4425/B sky130_fd_sc_hd__conb_1
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_831__883 VGND VGND VPWR VPWR _831__883/HI U$$4507/B sky130_fd_sc_hd__conb_1
XFILLER_48_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_52_2 dadda_fa_2_52_2/A dadda_fa_2_52_2/B dadda_fa_2_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/A dadda_fa_3_52_3/A sky130_fd_sc_hd__fa_2
XFILLER_39_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4040 U$$4040/A _675_/Q VGND VGND VPWR VPWR U$$4040/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_1 U$$2757/X U$$2890/X U$$3023/X VGND VGND VPWR VPWR dadda_fa_3_46_0/CIN
+ dadda_fa_3_45_2/CIN sky130_fd_sc_hd__fa_1
XU$$4051 U$$78/A1 U$$4107/A2 U$$765/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4052/A sky130_fd_sc_hd__a22o_1
XU$$4062 U$$4062/A _675_/Q VGND VGND VPWR VPWR U$$4062/X sky130_fd_sc_hd__xor2_1
XU$$4073 U$$4484/A1 U$$4107/A2 U$$4486/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4074/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4084 U$$4084/A U$$4109/A VGND VGND VPWR VPWR U$$4084/X sky130_fd_sc_hd__xor2_1
XU$$4095 U$$4506/A1 U$$4107/A2 U$$4508/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4096/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_0 dadda_fa_5_22_0/A dadda_fa_5_22_0/B dadda_fa_5_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/A dadda_fa_6_22_0/CIN sky130_fd_sc_hd__fa_1
XU$$3350 U$$3624/A1 U$$3412/A2 U$$3900/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3351/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_0 U$$1147/X U$$1280/X U$$1413/X VGND VGND VPWR VPWR dadda_fa_3_39_0/B
+ dadda_fa_3_38_2/B sky130_fd_sc_hd__fa_1
XU$$3361 U$$3361/A U$$3397/B VGND VGND VPWR VPWR U$$3361/X sky130_fd_sc_hd__xor2_1
XFILLER_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3372 U$$632/A1 U$$3412/A2 U$$771/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3373/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3383 U$$3383/A U$$3403/B VGND VGND VPWR VPWR U$$3383/X sky130_fd_sc_hd__xor2_1
XU$$3394 _601_/Q U$$3412/A2 U$$4492/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3395/A sky130_fd_sc_hd__a22o_1
XFILLER_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2660 U$$2660/A U$$2694/B VGND VGND VPWR VPWR U$$2660/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2671 U$$3217/B1 U$$2729/A2 U$$892/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2672/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2682 U$$2682/A U$$2698/B VGND VGND VPWR VPWR U$$2682/X sky130_fd_sc_hd__xor2_1
XU$$2693 U$$912/A1 U$$2729/A2 U$$914/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2694/A sky130_fd_sc_hd__a22o_1
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1970 U$$2790/B1 U$$2048/A2 U$$876/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1971/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1981 U$$1981/A U$$1991/B VGND VGND VPWR VPWR U$$1981/X sky130_fd_sc_hd__xor2_1
XU$$1992 U$$74/A1 U$$2048/A2 U$$76/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1993/A sky130_fd_sc_hd__a22o_1
XFILLER_21_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_67_2 dadda_fa_4_67_2/A dadda_fa_4_67_2/B dadda_fa_4_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/CIN dadda_fa_5_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput106 b[47] VGND VGND VPWR VPWR _599_/D sky130_fd_sc_hd__clkbuf_1
Xinput117 b[57] VGND VGND VPWR VPWR _609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput128 b[9] VGND VGND VPWR VPWR _561_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_193_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput139 c[109] VGND VGND VPWR VPWR input139/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$611 final_adder.U$$738/A final_adder.U$$738/B final_adder.U$$611/B1
+ VGND VGND VPWR VPWR final_adder.U$$739/B sky130_fd_sc_hd__a21o_1
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_37_0 dadda_fa_7_37_0/A dadda_fa_7_37_0/B dadda_fa_7_37_0/CIN VGND VGND
+ VPWR VPWR _462_/D _333_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$622 final_adder.U$$622/A _847__899/LO VGND VGND VPWR VPWR _168_/D
+ sky130_fd_sc_hd__xor2_2
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$633 final_adder.U$$633/A final_adder.U$$633/B VGND VGND VPWR VPWR
+ _179_/D sky130_fd_sc_hd__xor2_2
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$644 final_adder.U$$644/A final_adder.U$$644/B VGND VGND VPWR VPWR
+ _190_/D sky130_fd_sc_hd__xor2_2
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$655 final_adder.U$$655/A final_adder.U$$655/B VGND VGND VPWR VPWR
+ _201_/D sky130_fd_sc_hd__xor2_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$666 final_adder.U$$666/A final_adder.U$$666/B VGND VGND VPWR VPWR
+ _212_/D sky130_fd_sc_hd__xor2_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$505 U$$94/A1 U$$545/A2 U$$94/B1 U$$416/X VGND VGND VPWR VPWR U$$506/A sky130_fd_sc_hd__a22o_1
XFILLER_56_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$677 final_adder.U$$677/A final_adder.U$$677/B VGND VGND VPWR VPWR
+ _223_/D sky130_fd_sc_hd__xor2_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$516 U$$516/A U$$547/A VGND VGND VPWR VPWR U$$516/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_40_0 U$$87/X U$$220/X U$$353/X VGND VGND VPWR VPWR dadda_fa_2_41_3/CIN
+ dadda_fa_2_40_5/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$688 final_adder.U$$688/A final_adder.U$$688/B VGND VGND VPWR VPWR
+ _234_/D sky130_fd_sc_hd__xor2_1
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$527 U$$938/A1 U$$545/A2 U$$940/A1 U$$416/X VGND VGND VPWR VPWR U$$528/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$699 final_adder.U$$699/A final_adder.U$$699/B VGND VGND VPWR VPWR
+ _245_/D sky130_fd_sc_hd__xor2_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$538 U$$538/A _623_/Q VGND VGND VPWR VPWR U$$538/X sky130_fd_sc_hd__xor2_1
XU$$549 _624_/Q VGND VGND VPWR VPWR U$$551/B sky130_fd_sc_hd__inv_1
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_774__826 VGND VGND VPWR VPWR _774__826/HI U$$4393/B sky130_fd_sc_hd__conb_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_815__867 VGND VGND VPWR VPWR _815__867/HI U$$4475/B sky130_fd_sc_hd__conb_1
XFILLER_180_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_62_1 dadda_fa_3_62_1/A dadda_fa_3_62_1/B dadda_fa_3_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/CIN dadda_fa_4_62_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_55_0 dadda_fa_3_55_0/A dadda_fa_3_55_0/B dadda_fa_3_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/B dadda_fa_4_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1200 U$$787/B1 U$$1200/A2 U$$654/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1201/A sky130_fd_sc_hd__a22o_1
XFILLER_189_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1211 U$$1211/A U$$1232/A VGND VGND VPWR VPWR U$$1211/X sky130_fd_sc_hd__xor2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1222 U$$948/A1 U$$1100/X U$$950/A1 U$$1101/X VGND VGND VPWR VPWR U$$1223/A sky130_fd_sc_hd__a22o_1
XU$$1233 _633_/Q VGND VGND VPWR VPWR U$$1233/Y sky130_fd_sc_hd__inv_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1244 U$$1244/A U$$1336/B VGND VGND VPWR VPWR U$$1244/X sky130_fd_sc_hd__xor2_1
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1255 _559_/Q U$$1237/X U$$983/A1 U$$1238/X VGND VGND VPWR VPWR U$$1256/A sky130_fd_sc_hd__a22o_1
XU$$1266 U$$1266/A U$$1336/B VGND VGND VPWR VPWR U$$1266/X sky130_fd_sc_hd__xor2_1
XFILLER_31_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1277 U$$4291/A1 U$$1341/A2 U$$868/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1278/A
+ sky130_fd_sc_hd__a22o_1
XU$$1288 U$$1288/A U$$1336/B VGND VGND VPWR VPWR U$$1288/X sky130_fd_sc_hd__xor2_1
XU$$1299 U$$66/A1 U$$1341/A2 U$$68/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1300/A sky130_fd_sc_hd__a22o_1
XFILLER_176_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_112_0 dadda_fa_7_112_0/A dadda_fa_7_112_0/B dadda_fa_7_112_0/CIN VGND
+ VGND VPWR VPWR _537_/D _408_/D sky130_fd_sc_hd__fa_2
XFILLER_175_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_77_1 dadda_fa_5_77_1/A dadda_fa_5_77_1/B dadda_fa_5_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/B dadda_fa_7_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_8 dadda_fa_1_69_8/A dadda_fa_1_69_8/B dadda_fa_1_69_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_3/A dadda_fa_3_69_0/A sky130_fd_sc_hd__fa_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3180 U$$3180/A U$$3224/B VGND VGND VPWR VPWR U$$3180/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_9_0 dadda_fa_6_9_0/A dadda_fa_6_9_0/B dadda_fa_6_9_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_10_0/B dadda_fa_7_9_0/CIN sky130_fd_sc_hd__fa_2
XU$$3191 U$$3191/A1 U$$3241/A2 U$$3876/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3192/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2490 U$$4271/A1 U$$2534/A2 U$$4273/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_72_0 dadda_fa_4_72_0/A dadda_fa_4_72_0/B dadda_fa_4_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/A dadda_fa_5_72_1/A sky130_fd_sc_hd__fa_1
XFILLER_150_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_88_0 _689__909/HI U$$1779/X U$$1912/X VGND VGND VPWR VPWR dadda_fa_2_89_3/B
+ dadda_fa_2_88_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$441 final_adder.U$$264/B final_adder.U$$638/B final_adder.U$$145/X
+ VGND VGND VPWR VPWR final_adder.U$$640/B sky130_fd_sc_hd__a21o_1
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_621_ _621_/CLK _621_/D VGND VGND VPWR VPWR _621_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$463 final_adder.U$$286/B final_adder.U$$682/B final_adder.U$$189/X
+ VGND VGND VPWR VPWR final_adder.U$$684/B sky130_fd_sc_hd__a21o_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$302 U$$987/A1 U$$278/X U$$28/B1 U$$279/X VGND VGND VPWR VPWR U$$303/A sky130_fd_sc_hd__a22o_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$313 U$$313/A U$$391/B VGND VGND VPWR VPWR U$$313/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$485 final_adder.U$$308/B final_adder.U$$726/B final_adder.U$$233/X
+ VGND VGND VPWR VPWR final_adder.U$$728/B sky130_fd_sc_hd__a21o_1
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$324 U$$735/A1 U$$278/X U$$52/A1 U$$279/X VGND VGND VPWR VPWR U$$325/A sky130_fd_sc_hd__a22o_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$335 U$$335/A U$$357/B VGND VGND VPWR VPWR U$$335/X sky130_fd_sc_hd__xor2_1
X_552_ _576_/CLK _552_/D VGND VGND VPWR VPWR _552_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$346 U$$70/B1 U$$278/X U$$759/A1 U$$279/X VGND VGND VPWR VPWR U$$347/A sky130_fd_sc_hd__a22o_1
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$357 U$$357/A U$$357/B VGND VGND VPWR VPWR U$$357/X sky130_fd_sc_hd__xor2_1
XU$$368 U$$94/A1 U$$278/X U$$94/B1 U$$279/X VGND VGND VPWR VPWR U$$369/A sky130_fd_sc_hd__a22o_1
XFILLER_26_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$379 U$$379/A _621_/Q VGND VGND VPWR VPWR U$$379/X sky130_fd_sc_hd__xor2_1
XFILLER_83_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_483_ _483_/CLK _483_/D VGND VGND VPWR VPWR _483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_1_clk clkbuf_1_0_1_clk/A VGND VGND VPWR VPWR clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_87_0 dadda_fa_6_87_0/A dadda_fa_6_87_0/B dadda_fa_6_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_88_0/B dadda_fa_7_87_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_181_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$880 U$$880/A1 U$$910/A2 U$$60/A1 U$$910/B2 VGND VGND VPWR VPWR U$$881/A sky130_fd_sc_hd__a22o_1
XU$$1030 U$$1030/A U$$980/B VGND VGND VPWR VPWR U$$1030/X sky130_fd_sc_hd__xor2_1
XU$$891 U$$891/A U$$903/B VGND VGND VPWR VPWR U$$891/X sky130_fd_sc_hd__xor2_1
XU$$1041 U$$902/B1 U$$1093/A2 U$$84/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1042/A sky130_fd_sc_hd__a22o_1
XU$$1052 U$$1052/A U$$980/B VGND VGND VPWR VPWR U$$1052/X sky130_fd_sc_hd__xor2_1
XU$$1063 U$$787/B1 U$$1093/A2 U$$654/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1064/A sky130_fd_sc_hd__a22o_1
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1074 U$$1074/A _631_/Q VGND VGND VPWR VPWR U$$1074/X sky130_fd_sc_hd__xor2_1
XFILLER_177_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1085 U$$4510/A1 U$$1093/A2 _612_/Q U$$964/X VGND VGND VPWR VPWR U$$1086/A sky130_fd_sc_hd__a22o_1
XFILLER_188_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1096 U$$998/B VGND VGND VPWR VPWR U$$1096/Y sky130_fd_sc_hd__inv_1
XFILLER_192_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_81_7 U$$4026/X U$$4159/X U$$4292/X VGND VGND VPWR VPWR dadda_fa_2_82_3/B
+ dadda_fa_3_81_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_74_6 U$$4145/X U$$4278/X U$$4411/X VGND VGND VPWR VPWR dadda_fa_2_75_2/B
+ dadda_fa_2_74_5/B sky130_fd_sc_hd__fa_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_67_5 input220/X dadda_fa_1_67_5/B dadda_fa_1_67_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_68_2/A dadda_fa_2_67_5/A sky130_fd_sc_hd__fa_2
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_4 U$$1727/X U$$1860/X U$$1993/X VGND VGND VPWR VPWR dadda_fa_1_63_6/CIN
+ dadda_fa_1_62_8/CIN sky130_fd_sc_hd__fa_2
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3905 U$$3905/A U$$3929/B VGND VGND VPWR VPWR U$$3905/X sky130_fd_sc_hd__xor2_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_19_2 U$$843/X U$$976/X VGND VGND VPWR VPWR dadda_fa_4_20_1/B dadda_ha_3_19_2/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3916 U$$765/A1 U$$3970/A2 U$$82/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3917/A sky130_fd_sc_hd__a22o_1
XFILLER_40_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$260 final_adder.U$$260/A final_adder.U$$260/B VGND VGND VPWR VPWR
+ final_adder.U$$322/B sky130_fd_sc_hd__and2_1
XU$$3927 U$$3927/A _673_/Q VGND VGND VPWR VPWR U$$3927/X sky130_fd_sc_hd__xor2_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3938 U$$4486/A1 U$$3970/A2 U$$787/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3939/A
+ sky130_fd_sc_hd__a22o_1
XU$$110 _603_/Q U$$4/X U$$934/A1 U$$5/X VGND VGND VPWR VPWR U$$111/A sky130_fd_sc_hd__a22o_1
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_604_ _611_/CLK _604_/D VGND VGND VPWR VPWR _604_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$271 final_adder.U$$270/A final_adder.U$$157/X final_adder.U$$159/X
+ VGND VGND VPWR VPWR final_adder.U$$271/X sky130_fd_sc_hd__a21o_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3949 U$$3949/A U$$3969/B VGND VGND VPWR VPWR U$$3949/X sky130_fd_sc_hd__xor2_2
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$282 final_adder.U$$282/A final_adder.U$$282/B VGND VGND VPWR VPWR
+ final_adder.U$$332/A sky130_fd_sc_hd__and2_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_32_2 dadda_fa_3_32_2/A dadda_fa_3_32_2/B dadda_fa_3_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/A dadda_fa_4_32_2/B sky130_fd_sc_hd__fa_2
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$121 U$$121/A _617_/Q VGND VGND VPWR VPWR U$$121/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$293 final_adder.U$$292/A final_adder.U$$201/X final_adder.U$$203/X
+ VGND VGND VPWR VPWR final_adder.U$$293/X sky130_fd_sc_hd__a21o_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$132 U$$952/B1 U$$4/X U$$819/A1 U$$5/X VGND VGND VPWR VPWR U$$133/A sky130_fd_sc_hd__a22o_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$143 U$$143/A1 U$$141/X U$$8/A1 U$$142/X VGND VGND VPWR VPWR U$$144/A sky130_fd_sc_hd__a22o_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$154 U$$154/A U$$242/B VGND VGND VPWR VPWR U$$154/X sky130_fd_sc_hd__xor2_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_1 U$$1121/X U$$1254/X U$$1387/X VGND VGND VPWR VPWR dadda_fa_4_26_0/CIN
+ dadda_fa_4_25_2/A sky130_fd_sc_hd__fa_1
XFILLER_75_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_535_ _535_/CLK _535_/D VGND VGND VPWR VPWR _535_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$165 U$$28/A1 U$$141/X U$$28/B1 U$$142/X VGND VGND VPWR VPWR U$$166/A sky130_fd_sc_hd__a22o_1
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$176 U$$176/A U$$262/B VGND VGND VPWR VPWR U$$176/X sky130_fd_sc_hd__xor2_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$187 U$$735/A1 U$$141/X U$$52/A1 U$$142/X VGND VGND VPWR VPWR U$$188/A sky130_fd_sc_hd__a22o_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$198 U$$198/A U$$274/A VGND VGND VPWR VPWR U$$198/X sky130_fd_sc_hd__xor2_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_18_0 U$$43/X U$$176/X U$$309/X VGND VGND VPWR VPWR dadda_fa_4_19_1/A dadda_fa_4_18_2/A
+ sky130_fd_sc_hd__fa_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_466_ _467_/CLK _466_/D VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_397_ _535_/CLK _397_/D VGND VGND VPWR VPWR _397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_84_5 dadda_fa_2_84_5/A dadda_fa_2_84_5/B dadda_fa_2_84_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_2/A dadda_fa_4_84_0/A sky130_fd_sc_hd__fa_2
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_77_4 dadda_fa_2_77_4/A dadda_fa_2_77_4/B dadda_fa_2_77_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/CIN dadda_fa_3_77_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_100_3 U$$3665/X U$$3798/X U$$3931/X VGND VGND VPWR VPWR dadda_fa_3_101_2/B
+ dadda_fa_3_100_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_114_1 dadda_fa_5_114_1/A dadda_fa_5_114_1/B dadda_fa_5_114_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/B dadda_fa_7_114_0/A sky130_fd_sc_hd__fa_1
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_107_0 dadda_fa_5_107_0/A dadda_fa_5_107_0/B dadda_fa_5_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/A dadda_fa_6_107_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_133_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_72_3 U$$3210/X U$$3343/X U$$3476/X VGND VGND VPWR VPWR dadda_fa_2_73_1/B
+ dadda_fa_2_72_4/B sky130_fd_sc_hd__fa_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_65_2 U$$3329/X U$$3462/X U$$3595/X VGND VGND VPWR VPWR dadda_fa_2_66_1/A
+ dadda_fa_2_65_4/A sky130_fd_sc_hd__fa_1
XFILLER_87_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_42_1 dadda_fa_4_42_1/A dadda_fa_4_42_1/B dadda_fa_4_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/B dadda_fa_5_42_1/B sky130_fd_sc_hd__fa_1
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_58_1 U$$1985/X U$$2118/X U$$2251/X VGND VGND VPWR VPWR dadda_fa_2_59_0/CIN
+ dadda_fa_2_58_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_35_0 dadda_fa_4_35_0/A dadda_fa_4_35_0/B dadda_fa_4_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/A dadda_fa_5_35_1/A sky130_fd_sc_hd__fa_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_320_ _448_/CLK _320_/D VGND VGND VPWR VPWR _320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_251_ _503_/CLK _251_/D VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_182_ _458_/CLK hold4/X VGND VGND VPWR VPWR _182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_87_3 dadda_fa_3_87_3/A dadda_fa_3_87_3/B dadda_fa_3_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/B dadda_fa_4_87_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_136_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4403 U$$4403/A U$$4403/B VGND VGND VPWR VPWR U$$4403/X sky130_fd_sc_hd__xor2_2
XU$$4414 _563_/Q U$$4388/X _564_/Q U$$4389/X VGND VGND VPWR VPWR U$$4415/A sky130_fd_sc_hd__a22o_1
XU$$4425 U$$4425/A U$$4425/B VGND VGND VPWR VPWR U$$4425/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_60_1 U$$526/X U$$659/X U$$792/X VGND VGND VPWR VPWR dadda_fa_1_61_6/B
+ dadda_fa_1_60_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4436 _574_/Q U$$4388/X U$$4438/A1 U$$4389/X VGND VGND VPWR VPWR U$$4437/A sky130_fd_sc_hd__a22o_1
XU$$4447 U$$4447/A U$$4447/B VGND VGND VPWR VPWR U$$4447/X sky130_fd_sc_hd__xor2_1
XU$$3702 _671_/Q U$$3702/B VGND VGND VPWR VPWR U$$3702/X sky130_fd_sc_hd__and2_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4458 U$$759/A1 U$$4388/X U$$759/B1 U$$4389/X VGND VGND VPWR VPWR U$$4459/A sky130_fd_sc_hd__a22o_2
XU$$3713 U$$14/A1 U$$3783/A2 U$$14/B1 U$$3783/B2 VGND VGND VPWR VPWR U$$3714/A sky130_fd_sc_hd__a22o_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4469 U$$4469/A U$$4469/B VGND VGND VPWR VPWR U$$4469/X sky130_fd_sc_hd__xor2_2
XU$$3724 U$$3724/A U$$3756/B VGND VGND VPWR VPWR U$$3724/X sky130_fd_sc_hd__xor2_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3735 U$$4283/A1 U$$3783/A2 U$$4285/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3736/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3746 U$$3746/A U$$3784/B VGND VGND VPWR VPWR U$$3746/X sky130_fd_sc_hd__xor2_1
XFILLER_80_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3757 U$$4442/A1 U$$3795/A2 U$$4170/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3758/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_109_2 dadda_fa_4_109_2/A dadda_fa_4_109_2/B dadda_fa_4_109_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/CIN dadda_fa_5_109_1/CIN sky130_fd_sc_hd__fa_2
XU$$3768 U$$3768/A U$$3784/B VGND VGND VPWR VPWR U$$3768/X sky130_fd_sc_hd__xor2_1
XFILLER_79_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3779 _588_/Q U$$3795/A2 _589_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3780/A sky130_fd_sc_hd__a22o_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_518_ _518_/CLK _518_/D VGND VGND VPWR VPWR _518_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_449_ _461_/CLK _449_/D VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_82_2 dadda_fa_2_82_2/A dadda_fa_2_82_2/B dadda_fa_2_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/A dadda_fa_3_82_3/A sky130_fd_sc_hd__fa_1
XFILLER_173_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_75_1 dadda_fa_2_75_1/A dadda_fa_2_75_1/B dadda_fa_2_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/CIN dadda_fa_3_75_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_52_0 dadda_fa_5_52_0/A dadda_fa_5_52_0/B dadda_fa_5_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/A dadda_fa_6_52_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_123_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_68_0 dadda_fa_2_68_0/A dadda_fa_2_68_0/B dadda_fa_2_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/B dadda_fa_3_68_2/B sky130_fd_sc_hd__fa_2
XFILLER_29_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _367_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_97_2 dadda_fa_4_97_2/A dadda_fa_4_97_2/B dadda_fa_4_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/CIN dadda_fa_5_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_67_0 dadda_fa_7_67_0/A dadda_fa_7_67_0/B dadda_fa_7_67_0/CIN VGND VGND
+ VPWR VPWR _492_/D _363_/D sky130_fd_sc_hd__fa_2
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_70_0 U$$2275/X U$$2408/X U$$2541/X VGND VGND VPWR VPWR dadda_fa_2_71_0/B
+ dadda_fa_2_70_3/B sky130_fd_sc_hd__fa_2
XFILLER_120_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3009 U$$4379/A1 U$$3009/A2 U$$956/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$3010/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2308 _606_/Q U$$2316/A2 U$$940/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2309/A sky130_fd_sc_hd__a22o_1
XU$$2319 U$$2319/A U$$2327/B VGND VGND VPWR VPWR U$$2319/X sky130_fd_sc_hd__xor2_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1607 U$$98/B1 U$$1641/A2 U$$4486/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1608/A sky130_fd_sc_hd__a22o_1
XU$$1618 U$$1618/A U$$1643/A VGND VGND VPWR VPWR U$$1618/X sky130_fd_sc_hd__xor2_1
XU$$1629 U$$944/A1 U$$1641/A2 U$$946/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1630/A sky130_fd_sc_hd__a22o_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_742__794 VGND VGND VPWR VPWR _742__794/HI U$$2883/A1 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_81_clk _560_/CLK VGND VGND VPWR VPWR _637_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_303_ _303_/CLK _303_/D VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_234_ _499_/CLK _234_/D VGND VGND VPWR VPWR _234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_92_1 dadda_fa_3_92_1/A dadda_fa_3_92_1/B dadda_fa_3_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/CIN dadda_fa_4_92_2/A sky130_fd_sc_hd__fa_2
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_85_0 dadda_fa_3_85_0/A dadda_fa_3_85_0/B dadda_fa_3_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/B dadda_fa_4_85_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_136_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater507 U$$1512/X VGND VGND VPWR VPWR U$$1591/B2 sky130_fd_sc_hd__buf_12
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater518 U$$4247/A VGND VGND VPWR VPWR U$$4197/B sky130_fd_sc_hd__buf_12
XU$$4200 _593_/Q U$$4114/X U$$4476/A1 U$$4115/X VGND VGND VPWR VPWR U$$4201/A sky130_fd_sc_hd__a22o_1
Xrepeater529 _671_/Q VGND VGND VPWR VPWR U$$3794/B sky130_fd_sc_hd__buf_12
XFILLER_172_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4211 U$$4211/A _677_/Q VGND VGND VPWR VPWR U$$4211/X sky130_fd_sc_hd__xor2_1
XFILLER_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4222 U$$4496/A1 U$$4244/A2 U$$936/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4223/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4233 U$$4233/A U$$4246/A VGND VGND VPWR VPWR U$$4233/X sky130_fd_sc_hd__xor2_1
XU$$4244 U$$819/A1 U$$4244/A2 U$$4244/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4245/A
+ sky130_fd_sc_hd__a22o_1
XU$$3510 U$$3510/A U$$3536/B VGND VGND VPWR VPWR U$$3510/X sky130_fd_sc_hd__xor2_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_114_0 U$$4092/X U$$4225/X U$$4358/X VGND VGND VPWR VPWR dadda_fa_5_115_0/A
+ dadda_fa_5_114_1/A sky130_fd_sc_hd__fa_1
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_47_5 dadda_fa_2_47_5/A dadda_fa_2_47_5/B dadda_fa_2_47_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_2/A dadda_fa_4_47_0/A sky130_fd_sc_hd__fa_2
XU$$4255 U$$4255/A1 U$$4251/X _553_/Q U$$4252/X VGND VGND VPWR VPWR U$$4256/A sky130_fd_sc_hd__a22o_1
XU$$3521 _596_/Q U$$3545/A2 _597_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3522/A sky130_fd_sc_hd__a22o_1
XU$$4266 U$$4266/A U$$4332/B VGND VGND VPWR VPWR U$$4266/X sky130_fd_sc_hd__xor2_1
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4277 _563_/Q U$$4381/A2 _564_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4278/A sky130_fd_sc_hd__a22o_1
XU$$3532 U$$3532/A U$$3536/B VGND VGND VPWR VPWR U$$3532/X sky130_fd_sc_hd__xor2_1
XU$$4288 U$$4288/A U$$4384/A VGND VGND VPWR VPWR U$$4288/X sky130_fd_sc_hd__xor2_1
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3543 U$$4502/A1 U$$3429/X U$$4504/A1 U$$3430/X VGND VGND VPWR VPWR U$$3544/A sky130_fd_sc_hd__a22o_1
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3554 U$$3554/A U$$3561/A VGND VGND VPWR VPWR U$$3554/X sky130_fd_sc_hd__xor2_1
XU$$2820 _588_/Q U$$2870/A2 _589_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2821/A sky130_fd_sc_hd__a22o_1
XU$$4299 _574_/Q U$$4377/A2 U$$4438/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4300/A sky130_fd_sc_hd__a22o_1
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3565 _669_/Q U$$3565/B VGND VGND VPWR VPWR U$$3565/X sky130_fd_sc_hd__and2_1
XU$$3576 _555_/Q U$$3678/A2 U$$16/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3577/A sky130_fd_sc_hd__a22o_1
XU$$2831 U$$2831/A U$$2871/B VGND VGND VPWR VPWR U$$2831/X sky130_fd_sc_hd__xor2_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2842 _599_/Q U$$2868/A2 U$$926/A1 U$$2870/B2 VGND VGND VPWR VPWR U$$2843/A sky130_fd_sc_hd__a22o_1
XU$$3587 U$$3587/A U$$3625/B VGND VGND VPWR VPWR U$$3587/X sky130_fd_sc_hd__xor2_1
XFILLER_33_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3598 _566_/Q U$$3624/A2 _567_/Q U$$3624/B2 VGND VGND VPWR VPWR U$$3599/A sky130_fd_sc_hd__a22o_1
XU$$2853 U$$2853/A U$$2871/B VGND VGND VPWR VPWR U$$2853/X sky130_fd_sc_hd__xor2_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_clk _560_/CLK VGND VGND VPWR VPWR _579_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2864 _610_/Q U$$2870/A2 _611_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2865/A sky130_fd_sc_hd__a22o_1
XU$$2875 U$$2875/A _657_/Q VGND VGND VPWR VPWR U$$2875/X sky130_fd_sc_hd__xor2_1
XFILLER_178_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2886 U$$2886/A U$$2996/B VGND VGND VPWR VPWR U$$2886/X sky130_fd_sc_hd__xor2_1
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2897 U$$979/A1 U$$3009/A2 _559_/Q U$$3009/B2 VGND VGND VPWR VPWR U$$2898/A sky130_fd_sc_hd__a22o_1
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_691__911 VGND VGND VPWR VPWR _691__911/HI _691__911/LO sky130_fd_sc_hd__conb_1
XFILLER_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$709 _560_/Q U$$689/X U$$26/A1 U$$817/B2 VGND VGND VPWR VPWR U$$710/A sky130_fd_sc_hd__a22o_1
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_726__778 VGND VGND VPWR VPWR _726__778/HI U$$1924/A1 sky130_fd_sc_hd__conb_1
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _515_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_109_1 U$$3550/X U$$3683/X U$$3816/X VGND VGND VPWR VPWR dadda_fa_4_110_0/CIN
+ dadda_fa_4_109_2/A sky130_fd_sc_hd__fa_1
XFILLER_180_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2105 U$$50/A1 U$$2117/A2 U$$2790/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2106/A sky130_fd_sc_hd__a22o_1
XU$$2116 U$$2116/A U$$2118/B VGND VGND VPWR VPWR U$$2116/X sky130_fd_sc_hd__xor2_1
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2127 U$$70/B1 U$$2059/X U$$759/A1 U$$2060/X VGND VGND VPWR VPWR U$$2128/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2138 U$$2138/A _647_/Q VGND VGND VPWR VPWR U$$2138/X sky130_fd_sc_hd__xor2_1
XU$$2149 _595_/Q U$$2189/A2 _596_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2150/A sky130_fd_sc_hd__a22o_1
XU$$1404 U$$3457/B1 U$$1474/A2 U$$4283/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1405/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_54_clk _536_/CLK VGND VGND VPWR VPWR _537_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1415 U$$1415/A U$$1461/B VGND VGND VPWR VPWR U$$1415/X sky130_fd_sc_hd__xor2_1
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1426 U$$878/A1 U$$1472/A2 U$$880/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1427/A sky130_fd_sc_hd__a22o_1
XU$$1437 U$$1437/A U$$1479/B VGND VGND VPWR VPWR U$$1437/X sky130_fd_sc_hd__xor2_1
XU$$1448 U$$76/B1 U$$1472/A2 U$$902/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1449/A sky130_fd_sc_hd__a22o_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1459 U$$1459/A U$$1461/B VGND VGND VPWR VPWR U$$1459/X sky130_fd_sc_hd__xor2_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_217_ _480_/CLK _217_/D VGND VGND VPWR VPWR _217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_52_3 dadda_fa_2_52_3/A dadda_fa_2_52_3/B dadda_fa_2_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/B dadda_fa_3_52_3/B sky130_fd_sc_hd__fa_2
XU$$4030 U$$4030/A U$$4044/B VGND VGND VPWR VPWR U$$4030/X sky130_fd_sc_hd__xor2_1
XU$$4041 U$$4178/A1 U$$3977/X _583_/Q U$$3978/X VGND VGND VPWR VPWR U$$4042/A sky130_fd_sc_hd__a22o_1
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4052 U$$4052/A U$$4109/A VGND VGND VPWR VPWR U$$4052/X sky130_fd_sc_hd__xor2_1
XFILLER_38_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_45_2 input196/X dadda_fa_2_45_2/B dadda_fa_2_45_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_46_1/A dadda_fa_3_45_3/A sky130_fd_sc_hd__fa_2
XU$$4063 _593_/Q U$$4107/A2 U$$4476/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$4064/A sky130_fd_sc_hd__a22o_1
XU$$4074 U$$4074/A U$$4109/A VGND VGND VPWR VPWR U$$4074/X sky130_fd_sc_hd__xor2_1
XU$$3340 U$$50/B1 U$$3396/A2 U$$4438/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3341/A sky130_fd_sc_hd__a22o_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4085 U$$4496/A1 U$$4107/A2 _605_/Q U$$4107/B2 VGND VGND VPWR VPWR U$$4086/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_1 dadda_fa_5_22_1/A dadda_fa_5_22_1/B dadda_fa_5_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/B dadda_fa_7_22_0/A sky130_fd_sc_hd__fa_2
XU$$4096 U$$4096/A U$$4109/A VGND VGND VPWR VPWR U$$4096/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3351 U$$3351/A U$$3397/B VGND VGND VPWR VPWR U$$3351/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_38_1 U$$1546/X U$$1679/X U$$1812/X VGND VGND VPWR VPWR dadda_fa_3_39_0/CIN
+ dadda_fa_3_38_2/CIN sky130_fd_sc_hd__fa_2
XU$$3362 U$$4045/B1 U$$3396/A2 U$$76/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3363/A sky130_fd_sc_hd__a22o_1
XU$$3373 U$$3373/A U$$3413/B VGND VGND VPWR VPWR U$$3373/X sky130_fd_sc_hd__xor2_1
XU$$3384 U$$94/B1 U$$3412/A2 U$$98/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3385/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_45_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _280_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_5_15_0 dadda_fa_5_15_0/A dadda_fa_5_15_0/B dadda_fa_5_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/A dadda_fa_6_15_0/CIN sky130_fd_sc_hd__fa_1
XU$$2650 U$$2650/A U$$2698/B VGND VGND VPWR VPWR U$$2650/X sky130_fd_sc_hd__xor2_1
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3395 U$$3395/A U$$3413/B VGND VGND VPWR VPWR U$$3395/X sky130_fd_sc_hd__xor2_1
XFILLER_34_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2661 U$$58/A1 U$$2729/A2 _578_/Q U$$2729/B2 VGND VGND VPWR VPWR U$$2662/A sky130_fd_sc_hd__a22o_1
XFILLER_55_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2672 U$$2672/A U$$2694/B VGND VGND VPWR VPWR U$$2672/X sky130_fd_sc_hd__xor2_1
XU$$2683 U$$902/A1 U$$2729/A2 U$$902/B1 U$$2729/B2 VGND VGND VPWR VPWR U$$2684/A sky130_fd_sc_hd__a22o_1
XFILLER_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2694 U$$2694/A U$$2694/B VGND VGND VPWR VPWR U$$2694/X sky130_fd_sc_hd__xor2_1
XU$$1960 U$$3876/B1 U$$2048/A2 U$$4291/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1961/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1971 U$$1971/A U$$1991/B VGND VGND VPWR VPWR U$$1971/X sky130_fd_sc_hd__xor2_1
XU$$1982 U$$3900/A1 U$$2036/A2 U$$3489/B1 U$$2036/B2 VGND VGND VPWR VPWR U$$1983/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1993 U$$1993/A U$$2023/B VGND VGND VPWR VPWR U$$1993/X sky130_fd_sc_hd__xor2_1
XFILLER_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput107 b[48] VGND VGND VPWR VPWR _600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_41_3 U$$1286/X U$$1419/X VGND VGND VPWR VPWR dadda_fa_2_42_4/B dadda_fa_3_41_0/A
+ sky130_fd_sc_hd__ha_2
Xinput118 b[58] VGND VGND VPWR VPWR _610_/D sky130_fd_sc_hd__clkbuf_1
Xinput129 c[0] VGND VGND VPWR VPWR _424_/D sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$601 final_adder.U$$728/A final_adder.U$$728/B final_adder.U$$601/B1
+ VGND VGND VPWR VPWR final_adder.U$$729/B sky130_fd_sc_hd__a21o_1
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$623 final_adder.U$$623/A final_adder.U$$623/B VGND VGND VPWR VPWR
+ _169_/D sky130_fd_sc_hd__xor2_2
XFILLER_116_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$634 final_adder.U$$634/A final_adder.U$$634/B VGND VGND VPWR VPWR
+ _180_/D sky130_fd_sc_hd__xor2_1
Xdadda_ha_4_11_1 U$$428/X U$$561/X VGND VGND VPWR VPWR dadda_fa_5_12_0/CIN dadda_ha_4_11_1/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$645 final_adder.U$$645/A final_adder.U$$645/B VGND VGND VPWR VPWR
+ _191_/D sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$656 final_adder.U$$656/A final_adder.U$$656/B VGND VGND VPWR VPWR
+ _202_/D sky130_fd_sc_hd__xor2_1
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$667 final_adder.U$$667/A final_adder.U$$667/B VGND VGND VPWR VPWR
+ _213_/D sky130_fd_sc_hd__xor2_1
XFILLER_186_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$506 U$$506/A _623_/Q VGND VGND VPWR VPWR U$$506/X sky130_fd_sc_hd__xor2_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$678 final_adder.U$$678/A final_adder.U$$678/B VGND VGND VPWR VPWR
+ _224_/D sky130_fd_sc_hd__xor2_1
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$517 U$$928/A1 U$$545/A2 U$$930/A1 U$$416/X VGND VGND VPWR VPWR U$$518/A sky130_fd_sc_hd__a22o_1
XFILLER_84_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$689 final_adder.U$$689/A final_adder.U$$689/B VGND VGND VPWR VPWR
+ hold1/A sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_40_1 U$$486/X U$$619/X U$$752/X VGND VGND VPWR VPWR dadda_fa_2_41_4/A
+ dadda_fa_2_40_5/B sky130_fd_sc_hd__fa_2
XU$$528 U$$528/A U$$547/A VGND VGND VPWR VPWR U$$528/X sky130_fd_sc_hd__xor2_1
XU$$539 U$$539/A1 U$$415/X U$$952/A1 U$$416/X VGND VGND VPWR VPWR U$$540/A sky130_fd_sc_hd__a22o_1
XFILLER_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_clk _369_/CLK VGND VGND VPWR VPWR _499_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_62_2 dadda_fa_3_62_2/A dadda_fa_3_62_2/B dadda_fa_3_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/A dadda_fa_4_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_55_1 dadda_fa_3_55_1/A dadda_fa_3_55_1/B dadda_fa_3_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/CIN dadda_fa_4_55_2/A sky130_fd_sc_hd__fa_1
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_32_0 dadda_fa_6_32_0/A dadda_fa_6_32_0/B dadda_fa_6_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_33_0/B dadda_fa_7_32_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_48_0 dadda_fa_3_48_0/A dadda_fa_3_48_0/B dadda_fa_3_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/B dadda_fa_4_48_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk _369_/CLK VGND VGND VPWR VPWR _474_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1201 U$$1201/A _633_/Q VGND VGND VPWR VPWR U$$1201/X sky130_fd_sc_hd__xor2_1
XFILLER_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1212 _606_/Q U$$1100/X U$$940/A1 U$$1101/X VGND VGND VPWR VPWR U$$1213/A sky130_fd_sc_hd__a22o_1
XFILLER_189_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1223 U$$1223/A U$$1232/A VGND VGND VPWR VPWR U$$1223/X sky130_fd_sc_hd__xor2_1
XU$$1234 _634_/Q VGND VGND VPWR VPWR U$$1236/B sky130_fd_sc_hd__inv_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1245 U$$12/A1 U$$1341/A2 U$$14/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1246/A sky130_fd_sc_hd__a22o_1
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1256 U$$1256/A U$$1336/B VGND VGND VPWR VPWR U$$1256/X sky130_fd_sc_hd__xor2_1
XFILLER_149_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1267 U$$3457/B1 U$$1341/A2 U$$36/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1268/A sky130_fd_sc_hd__a22o_1
XFILLER_149_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1278 U$$1278/A U$$1342/B VGND VGND VPWR VPWR U$$1278/X sky130_fd_sc_hd__xor2_1
XFILLER_70_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1289 U$$878/A1 U$$1341/A2 U$$58/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1290/A sky130_fd_sc_hd__a22o_1
XFILLER_31_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_105_0 dadda_fa_7_105_0/A dadda_fa_7_105_0/B dadda_fa_7_105_0/CIN VGND
+ VGND VPWR VPWR _530_/D _401_/D sky130_fd_sc_hd__fa_2
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_0 U$$3496/B input202/X dadda_fa_2_50_0/CIN VGND VGND VPWR VPWR dadda_fa_3_51_0/B
+ dadda_fa_3_50_2/B sky130_fd_sc_hd__fa_2
XFILLER_39_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _462_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3170 U$$3170/A U$$3244/B VGND VGND VPWR VPWR U$$3170/X sky130_fd_sc_hd__xor2_1
XFILLER_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3181 _563_/Q U$$3243/A2 _564_/Q U$$3243/B2 VGND VGND VPWR VPWR U$$3182/A sky130_fd_sc_hd__a22o_1
XU$$3192 U$$3192/A U$$3224/B VGND VGND VPWR VPWR U$$3192/X sky130_fd_sc_hd__xor2_1
XFILLER_22_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_797__849 VGND VGND VPWR VPWR _797__849/HI U$$4439/B sky130_fd_sc_hd__conb_1
XFILLER_179_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2480 U$$12/B1 U$$2574/A2 U$$16/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2481/A sky130_fd_sc_hd__a22o_1
XU$$2491 U$$2491/A U$$2533/B VGND VGND VPWR VPWR U$$2491/X sky130_fd_sc_hd__xor2_1
XFILLER_50_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1790 U$$1790/A U$$1918/A VGND VGND VPWR VPWR U$$1790/X sky130_fd_sc_hd__xor2_1
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_72_1 dadda_fa_4_72_1/A dadda_fa_4_72_1/B dadda_fa_4_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/B dadda_fa_5_72_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_88_1 U$$2045/X U$$2178/X U$$2311/X VGND VGND VPWR VPWR dadda_fa_2_89_3/CIN
+ dadda_fa_2_88_5/A sky130_fd_sc_hd__fa_2
XFILLER_89_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_65_0 dadda_fa_4_65_0/A dadda_fa_4_65_0/B dadda_fa_4_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/A dadda_fa_5_65_1/A sky130_fd_sc_hd__fa_1
XFILLER_77_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$431 final_adder.U$$348/B final_adder.U$$734/B final_adder.U$$313/X
+ VGND VGND VPWR VPWR final_adder.U$$738/B sky130_fd_sc_hd__a21o_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ _620_/CLK _620_/D VGND VGND VPWR VPWR _620_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$453 final_adder.U$$276/B final_adder.U$$662/B final_adder.U$$169/X
+ VGND VGND VPWR VPWR final_adder.U$$664/B sky130_fd_sc_hd__a21o_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$303 U$$303/A U$$391/B VGND VGND VPWR VPWR U$$303/X sky130_fd_sc_hd__xor2_1
XFILLER_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$475 final_adder.U$$298/B final_adder.U$$706/B final_adder.U$$213/X
+ VGND VGND VPWR VPWR final_adder.U$$708/B sky130_fd_sc_hd__a21o_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$314 U$$40/A1 U$$278/X _569_/Q U$$279/X VGND VGND VPWR VPWR U$$315/A sky130_fd_sc_hd__a22o_1
XFILLER_123_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$325 U$$325/A U$$391/B VGND VGND VPWR VPWR U$$325/X sky130_fd_sc_hd__xor2_1
X_551_ _551_/CLK _551_/D VGND VGND VPWR VPWR _551_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater690 _582_/Q VGND VGND VPWR VPWR U$$3217/B1 sky130_fd_sc_hd__buf_12
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$497 final_adder.U$$624/A final_adder.U$$624/B final_adder.U$$497/B1
+ VGND VGND VPWR VPWR final_adder.U$$625/B sky130_fd_sc_hd__a21o_1
XU$$336 U$$62/A1 U$$278/X U$$64/A1 U$$279/X VGND VGND VPWR VPWR U$$337/A sky130_fd_sc_hd__a22o_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$347 U$$347/A U$$391/B VGND VGND VPWR VPWR U$$347/X sky130_fd_sc_hd__xor2_1
XU$$358 U$$84/A1 U$$278/X U$$86/A1 U$$279/X VGND VGND VPWR VPWR U$$359/A sky130_fd_sc_hd__a22o_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$369 U$$369/A U$$391/B VGND VGND VPWR VPWR U$$369/X sky130_fd_sc_hd__xor2_1
XFILLER_38_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_482_ _490_/CLK _482_/D VGND VGND VPWR VPWR _482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$870 U$$48/A1 U$$910/A2 U$$50/A1 U$$910/B2 VGND VGND VPWR VPWR U$$871/A sky130_fd_sc_hd__a22o_1
XU$$1020 U$$1020/A U$$998/B VGND VGND VPWR VPWR U$$1020/X sky130_fd_sc_hd__xor2_1
XU$$881 U$$881/A U$$903/B VGND VGND VPWR VPWR U$$881/X sky130_fd_sc_hd__xor2_1
XU$$1031 U$$72/A1 U$$999/A2 U$$74/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1032/A sky130_fd_sc_hd__a22o_1
XU$$892 U$$892/A1 U$$910/A2 U$$892/B1 U$$910/B2 VGND VGND VPWR VPWR U$$893/A sky130_fd_sc_hd__a22o_1
XU$$1042 U$$1042/A U$$980/B VGND VGND VPWR VPWR U$$1042/X sky130_fd_sc_hd__xor2_1
XU$$1053 U$$94/A1 U$$1093/A2 U$$94/B1 U$$1073/B2 VGND VGND VPWR VPWR U$$1054/A sky130_fd_sc_hd__a22o_1
XFILLER_177_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1064 U$$1064/A U$$998/B VGND VGND VPWR VPWR U$$1064/X sky130_fd_sc_hd__xor2_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1075 U$$938/A1 U$$963/X U$$940/A1 U$$964/X VGND VGND VPWR VPWR U$$1076/A sky130_fd_sc_hd__a22o_1
XU$$1086 U$$1086/A _631_/Q VGND VGND VPWR VPWR U$$1086/X sky130_fd_sc_hd__xor2_1
XFILLER_177_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1097 _632_/Q VGND VGND VPWR VPWR U$$1099/B sky130_fd_sc_hd__inv_1
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_82_0 dadda_fa_5_82_0/A dadda_fa_5_82_0/B dadda_fa_5_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/A dadda_fa_6_82_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_98_0 _697__917/HI U$$2464/X U$$2597/X VGND VGND VPWR VPWR dadda_fa_3_99_0/CIN
+ dadda_fa_3_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_172_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clk _431_/CLK VGND VGND VPWR VPWR _465_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_74_7 input228/X dadda_fa_1_74_7/B dadda_fa_1_74_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_75_2/CIN dadda_fa_2_74_5/CIN sky130_fd_sc_hd__fa_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_6 dadda_fa_1_67_6/A dadda_fa_1_67_6/B dadda_fa_1_67_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/B dadda_fa_2_67_5/B sky130_fd_sc_hd__fa_2
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_94_1 U$$2456/X U$$2589/X VGND VGND VPWR VPWR dadda_fa_2_95_5/CIN dadda_fa_3_94_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_183_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_97_0 dadda_fa_7_97_0/A dadda_fa_7_97_0/B dadda_fa_7_97_0/CIN VGND VGND
+ VPWR VPWR _522_/D _393_/D sky130_fd_sc_hd__fa_1
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_112_0 dadda_fa_6_112_0/A dadda_fa_6_112_0/B dadda_fa_6_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_113_0/B dadda_fa_7_112_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3906 U$$70/A1 U$$3912/A2 _584_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3907/A sky130_fd_sc_hd__a22o_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3917 U$$3917/A U$$3969/B VGND VGND VPWR VPWR U$$3917/X sky130_fd_sc_hd__xor2_1
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$250 final_adder.U$$745/A final_adder.U$$744/A VGND VGND VPWR VPWR
+ final_adder.U$$316/A sky130_fd_sc_hd__and2_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3928 U$$4476/A1 U$$3840/X _595_/Q U$$3841/X VGND VGND VPWR VPWR U$$3929/A sky130_fd_sc_hd__a22o_1
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_603_ _611_/CLK _603_/D VGND VGND VPWR VPWR _603_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$261 final_adder.U$$260/A final_adder.U$$137/X final_adder.U$$139/X
+ VGND VGND VPWR VPWR final_adder.U$$261/X sky130_fd_sc_hd__a21o_1
XU$$100 U$$98/B1 U$$4/X U$$924/A1 U$$5/X VGND VGND VPWR VPWR U$$101/A sky130_fd_sc_hd__a22o_1
XU$$3939 U$$3939/A _673_/Q VGND VGND VPWR VPWR U$$3939/X sky130_fd_sc_hd__xor2_1
XFILLER_85_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$272 final_adder.U$$272/A final_adder.U$$272/B VGND VGND VPWR VPWR
+ final_adder.U$$328/B sky130_fd_sc_hd__and2_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$111 U$$111/A _617_/Q VGND VGND VPWR VPWR U$$111/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$283 final_adder.U$$282/A final_adder.U$$181/X final_adder.U$$183/X
+ VGND VGND VPWR VPWR final_adder.U$$283/X sky130_fd_sc_hd__a21o_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$122 U$$944/A1 U$$4/X U$$946/A1 U$$5/X VGND VGND VPWR VPWR U$$123/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_32_3 dadda_fa_3_32_3/A dadda_fa_3_32_3/B dadda_fa_3_32_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/B dadda_fa_4_32_2/CIN sky130_fd_sc_hd__fa_2
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$294 final_adder.U$$294/A final_adder.U$$294/B VGND VGND VPWR VPWR
+ final_adder.U$$338/A sky130_fd_sc_hd__and2_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$133 U$$133/A U$$89/B VGND VGND VPWR VPWR U$$133/X sky130_fd_sc_hd__xor2_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$144 U$$144/A U$$242/B VGND VGND VPWR VPWR U$$144/X sky130_fd_sc_hd__xor2_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_534_ _535_/CLK _534_/D VGND VGND VPWR VPWR _534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$155 U$$975/B1 U$$141/X U$$842/A1 U$$142/X VGND VGND VPWR VPWR U$$156/A sky130_fd_sc_hd__a22o_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$166 U$$166/A U$$242/B VGND VGND VPWR VPWR U$$166/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_25_2 U$$1520/X U$$1653/X input174/X VGND VGND VPWR VPWR dadda_fa_4_26_1/A
+ dadda_fa_4_25_2/B sky130_fd_sc_hd__fa_2
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$177 U$$40/A1 U$$141/X _569_/Q U$$142/X VGND VGND VPWR VPWR U$$178/A sky130_fd_sc_hd__a22o_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$188 U$$188/A U$$262/B VGND VGND VPWR VPWR U$$188/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_18_1 U$$442/X U$$575/X U$$708/X VGND VGND VPWR VPWR dadda_fa_4_19_1/B
+ dadda_fa_4_18_2/B sky130_fd_sc_hd__fa_1
XU$$199 U$$62/A1 U$$141/X U$$64/A1 U$$142/X VGND VGND VPWR VPWR U$$200/A sky130_fd_sc_hd__a22o_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _465_/CLK _465_/D VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_396_ _543_/CLK _396_/D VGND VGND VPWR VPWR _396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_77_5 dadda_fa_2_77_5/A dadda_fa_2_77_5/B dadda_fa_2_77_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_2/A dadda_fa_4_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_107_1 dadda_fa_5_107_1/A dadda_fa_5_107_1/B dadda_fa_5_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/B dadda_fa_7_107_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_72_4 U$$3609/X U$$3742/X U$$3875/X VGND VGND VPWR VPWR dadda_fa_2_73_1/CIN
+ dadda_fa_2_72_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_65_3 U$$3728/X U$$3861/X U$$3994/X VGND VGND VPWR VPWR dadda_fa_2_66_1/B
+ dadda_fa_2_65_4/B sky130_fd_sc_hd__fa_1
XFILLER_87_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_42_2 dadda_fa_4_42_2/A dadda_fa_4_42_2/B dadda_fa_4_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/CIN dadda_fa_5_42_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_58_2 U$$2384/X U$$2517/X U$$2650/X VGND VGND VPWR VPWR dadda_fa_2_59_1/A
+ dadda_fa_2_58_4/A sky130_fd_sc_hd__fa_1
XFILLER_74_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_35_1 dadda_fa_4_35_1/A dadda_fa_4_35_1/B dadda_fa_4_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/B dadda_fa_5_35_1/B sky130_fd_sc_hd__fa_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_12_0 dadda_fa_7_12_0/A dadda_fa_7_12_0/B dadda_fa_7_12_0/CIN VGND VGND
+ VPWR VPWR _437_/D _308_/D sky130_fd_sc_hd__fa_2
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_28_0 dadda_fa_4_28_0/A dadda_fa_4_28_0/B dadda_fa_4_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/A dadda_fa_5_28_1/A sky130_fd_sc_hd__fa_2
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ _503_/CLK _250_/D VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_181_ _458_/CLK _181_/D VGND VGND VPWR VPWR _181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_61_4 U$$1725/X U$$1858/X VGND VGND VPWR VPWR dadda_fa_1_62_7/A dadda_fa_2_61_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4404 _558_/Q U$$4388/X _559_/Q U$$4389/X VGND VGND VPWR VPWR U$$4405/A sky130_fd_sc_hd__a22o_2
XFILLER_78_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4415 U$$4415/A U$$4415/B VGND VGND VPWR VPWR U$$4415/X sky130_fd_sc_hd__xor2_1
XU$$4426 _569_/Q U$$4388/X _570_/Q U$$4389/X VGND VGND VPWR VPWR U$$4427/A sky130_fd_sc_hd__a22o_1
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_60_2 U$$925/X U$$1058/X U$$1191/X VGND VGND VPWR VPWR dadda_fa_1_61_6/CIN
+ dadda_fa_1_60_8/B sky130_fd_sc_hd__fa_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4437 U$$4437/A U$$4437/B VGND VGND VPWR VPWR U$$4437/X sky130_fd_sc_hd__xor2_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3703 U$$3701/Y _670_/Q U$$3699/A U$$3702/X U$$3699/Y VGND VGND VPWR VPWR U$$3703/X
+ sky130_fd_sc_hd__a32o_4
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4448 _580_/Q U$$4388/X _581_/Q U$$4389/X VGND VGND VPWR VPWR U$$4449/A sky130_fd_sc_hd__a22o_1
XFILLER_93_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4459 U$$4459/A U$$4459/B VGND VGND VPWR VPWR U$$4459/X sky130_fd_sc_hd__xor2_4
XU$$3714 U$$3714/A U$$3756/B VGND VGND VPWR VPWR U$$3714/X sky130_fd_sc_hd__xor2_1
XFILLER_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3725 _561_/Q U$$3783/A2 _562_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3726/A sky130_fd_sc_hd__a22o_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3736 U$$3736/A U$$3756/B VGND VGND VPWR VPWR U$$3736/X sky130_fd_sc_hd__xor2_1
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3747 _572_/Q U$$3783/A2 U$$735/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3748/A sky130_fd_sc_hd__a22o_1
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_0 U$$1929/X U$$2062/X U$$2186/B VGND VGND VPWR VPWR dadda_fa_4_31_0/B
+ dadda_fa_4_30_1/CIN sky130_fd_sc_hd__fa_2
XU$$3758 U$$3758/A U$$3794/B VGND VGND VPWR VPWR U$$3758/X sky130_fd_sc_hd__xor2_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3769 U$$70/A1 U$$3783/A2 U$$70/B1 U$$3783/B2 VGND VGND VPWR VPWR U$$3770/A sky130_fd_sc_hd__a22o_1
XFILLER_166_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_517_ _527_/CLK _517_/D VGND VGND VPWR VPWR _517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _448_/CLK _448_/D VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_379_ _379_/CLK _379_/D VGND VGND VPWR VPWR _379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_82_3 dadda_fa_2_82_3/A dadda_fa_2_82_3/B dadda_fa_2_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/B dadda_fa_3_82_3/B sky130_fd_sc_hd__fa_2
Xdadda_fa_2_75_2 dadda_fa_2_75_2/A dadda_fa_2_75_2/B dadda_fa_2_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/A dadda_fa_3_75_3/A sky130_fd_sc_hd__fa_2
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_52_1 dadda_fa_5_52_1/A dadda_fa_5_52_1/B dadda_fa_5_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/B dadda_fa_7_52_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_68_1 dadda_fa_2_68_1/A dadda_fa_2_68_1/B dadda_fa_2_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/CIN dadda_fa_3_68_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_45_0 dadda_fa_5_45_0/A dadda_fa_5_45_0/B dadda_fa_5_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/A dadda_fa_6_45_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_70_1 U$$2674/X U$$2807/X U$$2940/X VGND VGND VPWR VPWR dadda_fa_2_71_0/CIN
+ dadda_fa_2_70_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_160_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_0 U$$2394/X U$$2527/X U$$2660/X VGND VGND VPWR VPWR dadda_fa_2_64_0/B
+ dadda_fa_2_63_3/B sky130_fd_sc_hd__fa_2
XFILLER_75_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2309 U$$2309/A _649_/Q VGND VGND VPWR VPWR U$$2309/X sky130_fd_sc_hd__xor2_1
XFILLER_28_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1608 U$$1608/A U$$1614/B VGND VGND VPWR VPWR U$$1608/X sky130_fd_sc_hd__xor2_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1619 U$$4496/A1 U$$1641/A2 U$$799/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1620/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_302_ _429_/CLK _302_/D VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_233_ _499_/CLK _233_/D VGND VGND VPWR VPWR _233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_92_2 dadda_fa_3_92_2/A dadda_fa_3_92_2/B dadda_fa_3_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/A dadda_fa_4_92_2/B sky130_fd_sc_hd__fa_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_85_1 dadda_fa_3_85_1/A dadda_fa_3_85_1/B dadda_fa_3_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/CIN dadda_fa_4_85_2/A sky130_fd_sc_hd__fa_1
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_62_0 dadda_fa_6_62_0/A dadda_fa_6_62_0/B dadda_fa_6_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_63_0/B dadda_fa_7_62_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_123_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_78_0 dadda_fa_3_78_0/A dadda_fa_3_78_0/B dadda_fa_3_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/B dadda_fa_4_78_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_123_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_52_0 U$$111/X U$$244/X VGND VGND VPWR VPWR dadda_fa_1_53_8/CIN dadda_fa_2_52_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_105_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater508 U$$1512/X VGND VGND VPWR VPWR U$$1641/B2 sky130_fd_sc_hd__buf_12
XU$$4201 U$$4201/A _677_/Q VGND VGND VPWR VPWR U$$4201/X sky130_fd_sc_hd__xor2_1
Xrepeater519 _677_/Q VGND VGND VPWR VPWR U$$4247/A sky130_fd_sc_hd__buf_12
XU$$4212 U$$4486/A1 U$$4244/A2 U$$787/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4213/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4223 U$$4223/A _677_/Q VGND VGND VPWR VPWR U$$4223/X sky130_fd_sc_hd__xor2_1
XU$$4234 U$$4508/A1 U$$4244/A2 U$$4510/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4235/A
+ sky130_fd_sc_hd__a22o_1
XU$$3500 U$$3500/A U$$3536/B VGND VGND VPWR VPWR U$$3500/X sky130_fd_sc_hd__xor2_1
XU$$4245 U$$4245/A U$$4246/A VGND VGND VPWR VPWR U$$4245/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3511 _591_/Q U$$3545/A2 U$$4335/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3512/A sky130_fd_sc_hd__a22o_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4256 U$$4256/A U$$4332/B VGND VGND VPWR VPWR U$$4256/X sky130_fd_sc_hd__xor2_1
XU$$3522 U$$3522/A U$$3536/B VGND VGND VPWR VPWR U$$3522/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_114_1 U$$4491/X input145/X dadda_fa_4_114_1/CIN VGND VGND VPWR VPWR dadda_fa_5_115_0/B
+ dadda_fa_5_114_1/B sky130_fd_sc_hd__fa_1
XFILLER_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4267 U$$979/A1 U$$4251/X U$$22/A1 U$$4252/X VGND VGND VPWR VPWR U$$4268/A sky130_fd_sc_hd__a22o_1
XFILLER_81_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4278 U$$4278/A _679_/Q VGND VGND VPWR VPWR U$$4278/X sky130_fd_sc_hd__xor2_1
XFILLER_81_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3533 U$$928/B1 U$$3545/A2 U$$4494/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3534/A
+ sky130_fd_sc_hd__a22o_1
XU$$3544 U$$3544/A U$$3561/A VGND VGND VPWR VPWR U$$3544/X sky130_fd_sc_hd__xor2_1
XU$$4289 U$$4289/A1 U$$4251/X U$$4289/B1 U$$4252/X VGND VGND VPWR VPWR U$$4290/A sky130_fd_sc_hd__a22o_1
XU$$2810 _583_/Q U$$2870/A2 _584_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2811/A sky130_fd_sc_hd__a22o_1
XU$$3555 U$$4514/A1 U$$3429/X U$$4379/A1 U$$3430/X VGND VGND VPWR VPWR U$$3556/A sky130_fd_sc_hd__a22o_1
XU$$2821 U$$2821/A U$$2871/B VGND VGND VPWR VPWR U$$2821/X sky130_fd_sc_hd__xor2_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_107_0 dadda_fa_4_107_0/A dadda_fa_4_107_0/B dadda_fa_4_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/A dadda_fa_5_107_1/A sky130_fd_sc_hd__fa_2
XFILLER_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3566 U$$3564/Y _668_/Q _667_/Q U$$3565/X U$$3562/Y VGND VGND VPWR VPWR U$$3566/X
+ sky130_fd_sc_hd__a32o_4
XU$$2832 _594_/Q U$$2870/A2 _595_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2833/A sky130_fd_sc_hd__a22o_1
XU$$3577 U$$3577/A U$$3698/A VGND VGND VPWR VPWR U$$3577/X sky130_fd_sc_hd__xor2_1
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2843 U$$2843/A U$$2871/B VGND VGND VPWR VPWR U$$2843/X sky130_fd_sc_hd__xor2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3588 U$$4273/A1 U$$3624/A2 U$$28/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3589/A sky130_fd_sc_hd__a22o_1
XU$$2854 U$$936/A1 U$$2744/X _606_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2855/A sky130_fd_sc_hd__a22o_1
XFILLER_73_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3599 U$$3599/A U$$3625/B VGND VGND VPWR VPWR U$$3599/X sky130_fd_sc_hd__xor2_1
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2865 U$$2865/A U$$2871/B VGND VGND VPWR VPWR U$$2865/X sky130_fd_sc_hd__xor2_1
XFILLER_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2876 _657_/Q VGND VGND VPWR VPWR U$$2876/Y sky130_fd_sc_hd__inv_1
XU$$2887 _553_/Q U$$2975/A2 U$$4122/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2888/A sky130_fd_sc_hd__a22o_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2898 U$$2898/A U$$2996/B VGND VGND VPWR VPWR U$$2898/X sky130_fd_sc_hd__xor2_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_80_0 input235/X dadda_fa_2_80_0/B dadda_fa_2_80_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_81_0/B dadda_fa_3_80_2/B sky130_fd_sc_hd__fa_2
XFILLER_143_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_1_50_8 U$$3299/X U$$3432/X VGND VGND VPWR VPWR dadda_fa_2_51_3/A dadda_fa_3_50_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_95_0 dadda_fa_4_95_0/A dadda_fa_4_95_0/B dadda_fa_4_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/A dadda_fa_5_95_1/A sky130_fd_sc_hd__fa_2
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_109_2 U$$3949/X U$$4082/X U$$4215/X VGND VGND VPWR VPWR dadda_fa_4_110_1/A
+ dadda_fa_4_109_2/B sky130_fd_sc_hd__fa_2
XFILLER_180_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput380 _264_/Q VGND VGND VPWR VPWR o[96] sky130_fd_sc_hd__buf_2
XFILLER_160_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2106 U$$2106/A U$$2118/B VGND VGND VPWR VPWR U$$2106/X sky130_fd_sc_hd__xor2_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2117 U$$3624/A1 U$$2117/A2 U$$3900/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2118/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2128 U$$2128/A U$$2186/B VGND VGND VPWR VPWR U$$2128/X sky130_fd_sc_hd__xor2_1
XFILLER_16_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2139 U$$632/A1 U$$2161/A2 U$$771/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2140/A sky130_fd_sc_hd__a22o_1
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1405 U$$1405/A U$$1461/B VGND VGND VPWR VPWR U$$1405/X sky130_fd_sc_hd__xor2_1
XFILLER_55_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1416 U$$868/A1 U$$1472/A2 U$$48/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1417/A sky130_fd_sc_hd__a22o_1
XFILLER_167_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1427 U$$1427/A U$$1505/B VGND VGND VPWR VPWR U$$1427/X sky130_fd_sc_hd__xor2_1
XU$$1438 U$$3217/B1 U$$1472/A2 U$$892/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1439/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1449 U$$1449/A U$$1505/B VGND VGND VPWR VPWR U$$1449/X sky130_fd_sc_hd__xor2_1
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_216_ _456_/CLK _216_/D VGND VGND VPWR VPWR _216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_52_4 dadda_fa_2_52_4/A dadda_fa_2_52_4/B dadda_fa_2_52_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/CIN dadda_fa_3_52_3/CIN sky130_fd_sc_hd__fa_2
XU$$4020 U$$4020/A U$$4058/B VGND VGND VPWR VPWR U$$4020/X sky130_fd_sc_hd__xor2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4031 U$$4442/A1 U$$4045/A2 _578_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$4032/A sky130_fd_sc_hd__a22o_1
XU$$4042 U$$4042/A U$$4058/B VGND VGND VPWR VPWR U$$4042/X sky130_fd_sc_hd__xor2_1
XU$$4053 U$$765/A1 U$$3977/X _589_/Q U$$3978/X VGND VGND VPWR VPWR U$$4054/A sky130_fd_sc_hd__a22o_1
XFILLER_65_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_45_3 dadda_fa_2_45_3/A dadda_fa_2_45_3/B dadda_fa_2_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/B dadda_fa_3_45_3/B sky130_fd_sc_hd__fa_2
XU$$4064 U$$4064/A _675_/Q VGND VGND VPWR VPWR U$$4064/X sky130_fd_sc_hd__xor2_1
XU$$4075 U$$4486/A1 U$$4107/A2 U$$787/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4076/A
+ sky130_fd_sc_hd__a22o_1
XU$$3330 U$$4289/A1 U$$3412/A2 U$$4291/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3331/A
+ sky130_fd_sc_hd__a22o_1
XU$$3341 U$$3341/A U$$3397/B VGND VGND VPWR VPWR U$$3341/X sky130_fd_sc_hd__xor2_1
XU$$4086 U$$4086/A U$$4109/A VGND VGND VPWR VPWR U$$4086/X sky130_fd_sc_hd__xor2_1
XU$$3352 _580_/Q U$$3292/X _581_/Q U$$3293/X VGND VGND VPWR VPWR U$$3353/A sky130_fd_sc_hd__a22o_1
XU$$4097 U$$4508/A1 U$$4107/A2 U$$4510/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4098/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_2 U$$1945/X U$$2078/X U$$2211/X VGND VGND VPWR VPWR dadda_fa_3_39_1/A
+ dadda_fa_3_38_3/A sky130_fd_sc_hd__fa_2
XU$$3363 U$$3363/A U$$3397/B VGND VGND VPWR VPWR U$$3363/X sky130_fd_sc_hd__xor2_1
XU$$3374 U$$771/A1 U$$3412/A2 U$$771/B1 U$$3412/B2 VGND VGND VPWR VPWR U$$3375/A sky130_fd_sc_hd__a22o_1
XU$$2640 U$$2640/A U$$2694/B VGND VGND VPWR VPWR U$$2640/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_15_1 dadda_fa_5_15_1/A dadda_fa_5_15_1/B dadda_fa_5_15_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/B dadda_fa_7_15_0/A sky130_fd_sc_hd__fa_2
XU$$3385 U$$3385/A U$$3413/B VGND VGND VPWR VPWR U$$3385/X sky130_fd_sc_hd__xor2_1
XU$$2651 U$$4156/B1 U$$2607/X _573_/Q U$$2608/X VGND VGND VPWR VPWR U$$2652/A sky130_fd_sc_hd__a22o_1
XFILLER_0_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3396 U$$928/B1 U$$3396/A2 U$$4494/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3397/A
+ sky130_fd_sc_hd__a22o_1
XU$$2662 U$$2662/A U$$2710/B VGND VGND VPWR VPWR U$$2662/X sky130_fd_sc_hd__xor2_1
XFILLER_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2673 _583_/Q U$$2607/X _584_/Q U$$2608/X VGND VGND VPWR VPWR U$$2674/A sky130_fd_sc_hd__a22o_1
XU$$2684 U$$2684/A U$$2694/B VGND VGND VPWR VPWR U$$2684/X sky130_fd_sc_hd__xor2_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1950 U$$30/B1 U$$2048/A2 U$$3457/B1 U$$2048/B2 VGND VGND VPWR VPWR U$$1951/A sky130_fd_sc_hd__a22o_1
XU$$2695 U$$914/A1 U$$2729/A2 U$$92/B1 U$$2729/B2 VGND VGND VPWR VPWR U$$2696/A sky130_fd_sc_hd__a22o_1
XFILLER_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1961 U$$1961/A U$$1991/B VGND VGND VPWR VPWR U$$1961/X sky130_fd_sc_hd__xor2_1
XU$$1972 U$$4438/A1 U$$2036/A2 U$$878/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1973/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1983 U$$1983/A U$$1991/B VGND VGND VPWR VPWR U$$1983/X sky130_fd_sc_hd__xor2_1
XFILLER_22_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1994 U$$759/B1 U$$2048/A2 U$$78/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1995/A sky130_fd_sc_hd__a22o_1
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput108 b[49] VGND VGND VPWR VPWR _601_/D sky130_fd_sc_hd__clkbuf_1
Xinput119 b[59] VGND VGND VPWR VPWR _611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$613 final_adder.U$$740/A final_adder.U$$740/B final_adder.U$$613/B1
+ VGND VGND VPWR VPWR final_adder.U$$741/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$624 final_adder.U$$624/A final_adder.U$$624/B VGND VGND VPWR VPWR
+ _170_/D sky130_fd_sc_hd__xor2_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$635 final_adder.U$$635/A final_adder.U$$635/B VGND VGND VPWR VPWR
+ _181_/D sky130_fd_sc_hd__xor2_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$646 final_adder.U$$646/A final_adder.U$$646/B VGND VGND VPWR VPWR
+ _192_/D sky130_fd_sc_hd__xor2_1
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$657 final_adder.U$$657/A final_adder.U$$657/B VGND VGND VPWR VPWR
+ _203_/D sky130_fd_sc_hd__xor2_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$668 final_adder.U$$668/A final_adder.U$$668/B VGND VGND VPWR VPWR
+ _214_/D sky130_fd_sc_hd__xor2_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$507 U$$96/A1 U$$545/A2 U$$96/B1 U$$416/X VGND VGND VPWR VPWR U$$508/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$679 final_adder.U$$679/A final_adder.U$$679/B VGND VGND VPWR VPWR
+ _225_/D sky130_fd_sc_hd__xor2_1
XU$$518 U$$518/A U$$530/B VGND VGND VPWR VPWR U$$518/X sky130_fd_sc_hd__xor2_1
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$529 U$$940/A1 U$$545/A2 U$$942/A1 U$$416/X VGND VGND VPWR VPWR U$$530/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_40_2 U$$885/X U$$1018/X U$$1151/X VGND VGND VPWR VPWR dadda_fa_2_41_4/B
+ dadda_fa_2_40_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_698__918 VGND VGND VPWR VPWR _698__918/HI _698__918/LO sky130_fd_sc_hd__conb_1
XU$$90 U$$90/A1 U$$4/X U$$92/A1 U$$5/X VGND VGND VPWR VPWR U$$91/A sky130_fd_sc_hd__a22o_1
XFILLER_53_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_10_0 U$$27/X U$$160/X U$$293/X VGND VGND VPWR VPWR dadda_fa_5_11_0/CIN
+ dadda_fa_5_10_1/B sky130_fd_sc_hd__fa_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_114_0 _700__920/HI U$$3560/X U$$3693/X VGND VGND VPWR VPWR dadda_fa_4_115_2/A
+ dadda_fa_4_114_2/B sky130_fd_sc_hd__fa_1
XFILLER_119_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_62_3 dadda_fa_3_62_3/A dadda_fa_3_62_3/B dadda_fa_3_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/B dadda_fa_4_62_2/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_55_2 dadda_fa_3_55_2/A dadda_fa_3_55_2/B dadda_fa_3_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/A dadda_fa_4_55_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_3_48_1 dadda_fa_3_48_1/A dadda_fa_3_48_1/B dadda_fa_3_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/CIN dadda_fa_4_48_2/A sky130_fd_sc_hd__fa_1
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_25_0 dadda_fa_6_25_0/A dadda_fa_6_25_0/B dadda_fa_6_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_26_0/B dadda_fa_7_25_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_63_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1202 U$$654/A1 U$$1100/X U$$930/A1 U$$1101/X VGND VGND VPWR VPWR U$$1203/A sky130_fd_sc_hd__a22o_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1213 U$$1213/A U$$1232/A VGND VGND VPWR VPWR U$$1213/X sky130_fd_sc_hd__xor2_1
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1224 U$$539/A1 U$$1100/X U$$4514/A1 U$$1101/X VGND VGND VPWR VPWR U$$1225/A sky130_fd_sc_hd__a22o_1
XFILLER_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1235 _635_/Q VGND VGND VPWR VPWR U$$1235/Y sky130_fd_sc_hd__inv_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1246 U$$1246/A U$$1342/B VGND VGND VPWR VPWR U$$1246/X sky130_fd_sc_hd__xor2_1
XFILLER_31_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1257 U$$983/A1 U$$1237/X U$$26/A1 U$$1238/X VGND VGND VPWR VPWR U$$1258/A sky130_fd_sc_hd__a22o_1
XFILLER_43_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1268 U$$1268/A U$$1342/B VGND VGND VPWR VPWR U$$1268/X sky130_fd_sc_hd__xor2_1
XFILLER_176_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1279 U$$868/A1 U$$1341/A2 U$$48/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1280/A sky130_fd_sc_hd__a22o_1
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_1 dadda_fa_2_50_1/A dadda_fa_2_50_1/B dadda_fa_2_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_0/CIN dadda_fa_3_50_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_22_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_43_0 U$$1955/X U$$2088/X U$$2221/X VGND VGND VPWR VPWR dadda_fa_3_44_0/B
+ dadda_fa_3_43_2/B sky130_fd_sc_hd__fa_2
XFILLER_4_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3160 U$$3160/A U$$3224/B VGND VGND VPWR VPWR U$$3160/X sky130_fd_sc_hd__xor2_1
XU$$3171 U$$979/A1 U$$3243/A2 U$$979/B1 U$$3243/B2 VGND VGND VPWR VPWR U$$3172/A sky130_fd_sc_hd__a22o_1
XFILLER_179_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3182 U$$3182/A U$$3244/B VGND VGND VPWR VPWR U$$3182/X sky130_fd_sc_hd__xor2_1
XFILLER_35_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3193 U$$3876/B1 U$$3241/A2 U$$4291/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3194/A
+ sky130_fd_sc_hd__a22o_1
XU$$2470 U$$2468/Y _652_/Q _651_/Q U$$2469/X U$$2466/Y VGND VGND VPWR VPWR U$$2470/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2481 U$$2481/A U$$2533/B VGND VGND VPWR VPWR U$$2481/X sky130_fd_sc_hd__xor2_1
XFILLER_179_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2492 U$$4273/A1 U$$2534/A2 U$$28/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2493/A sky130_fd_sc_hd__a22o_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1780 _641_/Q VGND VGND VPWR VPWR U$$1780/Y sky130_fd_sc_hd__inv_1
XFILLER_107_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1791 U$$8/B1 U$$1867/A2 U$$971/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1792/A sky130_fd_sc_hd__a22o_1
XFILLER_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput90 b[32] VGND VGND VPWR VPWR _584_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_72_2 dadda_fa_4_72_2/A dadda_fa_4_72_2/B dadda_fa_4_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/CIN dadda_fa_5_72_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_88_2 U$$2444/X U$$2577/X U$$2710/X VGND VGND VPWR VPWR dadda_fa_2_89_4/A
+ dadda_fa_2_88_5/B sky130_fd_sc_hd__fa_1
XFILLER_27_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_65_1 dadda_fa_4_65_1/A dadda_fa_4_65_1/B dadda_fa_4_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/B dadda_fa_5_65_1/B sky130_fd_sc_hd__fa_1
XFILLER_104_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_42_0 dadda_fa_7_42_0/A dadda_fa_7_42_0/B dadda_fa_7_42_0/CIN VGND VGND
+ VPWR VPWR _467_/D _338_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_58_0 dadda_fa_4_58_0/A dadda_fa_4_58_0/B dadda_fa_4_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/A dadda_fa_5_58_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$421 final_adder.U$$338/B final_adder.U$$694/B final_adder.U$$293/X
+ VGND VGND VPWR VPWR final_adder.U$$698/B sky130_fd_sc_hd__a21o_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$443 final_adder.U$$266/B final_adder.U$$642/B final_adder.U$$149/X
+ VGND VGND VPWR VPWR final_adder.U$$644/B sky130_fd_sc_hd__a21o_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_780__832 VGND VGND VPWR VPWR _780__832/HI U$$4405/B sky130_fd_sc_hd__conb_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$465 final_adder.U$$288/B final_adder.U$$686/B final_adder.U$$193/X
+ VGND VGND VPWR VPWR final_adder.U$$688/B sky130_fd_sc_hd__a21o_1
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$304 U$$28/B1 U$$278/X U$$32/A1 U$$279/X VGND VGND VPWR VPWR U$$305/A sky130_fd_sc_hd__a22o_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_550_ _650_/CLK _550_/D VGND VGND VPWR VPWR _550_/Q sky130_fd_sc_hd__dfxtp_4
XU$$315 U$$315/A U$$357/B VGND VGND VPWR VPWR U$$315/X sky130_fd_sc_hd__xor2_1
Xrepeater680 U$$4045/B1 VGND VGND VPWR VPWR U$$74/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$487 final_adder.U$$310/B final_adder.U$$730/B final_adder.U$$237/X
+ VGND VGND VPWR VPWR final_adder.U$$732/B sky130_fd_sc_hd__a21o_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$326 U$$52/A1 U$$278/X U$$54/A1 U$$279/X VGND VGND VPWR VPWR U$$327/A sky130_fd_sc_hd__a22o_1
Xrepeater691 _582_/Q VGND VGND VPWR VPWR U$$4178/A1 sky130_fd_sc_hd__buf_12
XFILLER_123_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$337 U$$337/A U$$391/B VGND VGND VPWR VPWR U$$337/X sky130_fd_sc_hd__xor2_1
XFILLER_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$348 U$$759/A1 U$$278/X U$$759/B1 U$$279/X VGND VGND VPWR VPWR U$$349/A sky130_fd_sc_hd__a22o_1
XU$$359 U$$359/A U$$391/B VGND VGND VPWR VPWR U$$359/X sky130_fd_sc_hd__xor2_1
X_481_ _490_/CLK _481_/D VGND VGND VPWR VPWR _481_/Q sky130_fd_sc_hd__dfxtp_1
X_821__873 VGND VGND VPWR VPWR _821__873/HI U$$4487/B sky130_fd_sc_hd__conb_1
XFILLER_38_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_60_0 dadda_fa_3_60_0/A dadda_fa_3_60_0/B dadda_fa_3_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/B dadda_fa_4_60_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_76_0 _684__904/HI U$$957/X U$$1090/X VGND VGND VPWR VPWR dadda_fa_1_77_8/B
+ dadda_fa_1_76_8/CIN sky130_fd_sc_hd__fa_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$860 U$$38/A1 U$$928/A2 U$$40/A1 U$$928/B2 VGND VGND VPWR VPWR U$$861/A sky130_fd_sc_hd__a22o_1
XFILLER_17_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_679_ _679_/CLK _679_/D VGND VGND VPWR VPWR _679_/Q sky130_fd_sc_hd__dfxtp_4
XU$$1010 U$$1010/A U$$980/B VGND VGND VPWR VPWR U$$1010/X sky130_fd_sc_hd__xor2_1
XU$$871 U$$871/A U$$943/B VGND VGND VPWR VPWR U$$871/X sky130_fd_sc_hd__xor2_1
XFILLER_17_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1021 U$$62/A1 U$$999/A2 U$$64/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1022/A sky130_fd_sc_hd__a22o_1
XFILLER_16_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$882 U$$60/A1 U$$910/A2 U$$62/A1 U$$910/B2 VGND VGND VPWR VPWR U$$883/A sky130_fd_sc_hd__a22o_1
XFILLER_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1032 U$$1032/A U$$980/B VGND VGND VPWR VPWR U$$1032/X sky130_fd_sc_hd__xor2_1
XU$$893 U$$893/A U$$943/B VGND VGND VPWR VPWR U$$893/X sky130_fd_sc_hd__xor2_1
XFILLER_32_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1043 U$$84/A1 U$$999/A2 U$$86/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1044/A sky130_fd_sc_hd__a22o_1
XU$$1054 U$$1054/A U$$998/B VGND VGND VPWR VPWR U$$1054/X sky130_fd_sc_hd__xor2_1
XU$$1065 U$$654/A1 U$$963/X U$$930/A1 U$$964/X VGND VGND VPWR VPWR U$$1066/A sky130_fd_sc_hd__a22o_1
XFILLER_177_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1076 U$$1076/A _631_/Q VGND VGND VPWR VPWR U$$1076/X sky130_fd_sc_hd__xor2_1
XFILLER_189_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1087 _612_/Q U$$963/X U$$4514/A1 U$$964/X VGND VGND VPWR VPWR U$$1088/A sky130_fd_sc_hd__a22o_1
XU$$1098 _633_/Q VGND VGND VPWR VPWR U$$1098/Y sky130_fd_sc_hd__inv_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_82_1 dadda_fa_5_82_1/A dadda_fa_5_82_1/B dadda_fa_5_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/B dadda_fa_7_82_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_98_1 U$$2730/X U$$2863/X U$$2996/X VGND VGND VPWR VPWR dadda_fa_3_99_1/A
+ dadda_fa_3_98_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_75_0 dadda_fa_5_75_0/A dadda_fa_5_75_0/B dadda_fa_5_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/A dadda_fa_6_75_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_74_8 dadda_fa_1_74_8/A dadda_fa_1_74_8/B dadda_fa_1_74_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_75_3/A dadda_fa_3_74_0/A sky130_fd_sc_hd__fa_2
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_764__816 VGND VGND VPWR VPWR _764__816/HI U$$4244/B1 sky130_fd_sc_hd__conb_1
XFILLER_101_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_67_7 dadda_fa_1_67_7/A dadda_fa_1_67_7/B dadda_fa_1_67_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/CIN dadda_fa_2_67_5/CIN sky130_fd_sc_hd__fa_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_805__857 VGND VGND VPWR VPWR _805__857/HI U$$4455/B sky130_fd_sc_hd__conb_1
XFILLER_187_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_93_0 U$$2054/Y U$$2188/X U$$2321/X VGND VGND VPWR VPWR dadda_fa_2_94_5/A
+ dadda_fa_2_93_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3907 U$$3907/A U$$3929/B VGND VGND VPWR VPWR U$$3907/X sky130_fd_sc_hd__xor2_1
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$240 final_adder.U$$735/A final_adder.U$$734/A VGND VGND VPWR VPWR
+ final_adder.U$$312/B sky130_fd_sc_hd__and2_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$251 final_adder.U$$745/A final_adder.U$$617/B1 final_adder.U$$251/B1
+ VGND VGND VPWR VPWR final_adder.U$$251/X sky130_fd_sc_hd__a21o_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3918 U$$82/A1 U$$3970/A2 U$$632/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3919/A sky130_fd_sc_hd__a22o_1
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_602_ _611_/CLK _602_/D VGND VGND VPWR VPWR _602_/Q sky130_fd_sc_hd__dfxtp_4
XU$$101 U$$101/A U$$89/B VGND VGND VPWR VPWR U$$101/X sky130_fd_sc_hd__xor2_1
XFILLER_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3929 U$$3929/A U$$3929/B VGND VGND VPWR VPWR U$$3929/X sky130_fd_sc_hd__xor2_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$262 final_adder.U$$262/A final_adder.U$$262/B VGND VGND VPWR VPWR
+ final_adder.U$$322/A sky130_fd_sc_hd__and2_1
Xdadda_fa_6_105_0 dadda_fa_6_105_0/A dadda_fa_6_105_0/B dadda_fa_6_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_106_0/B dadda_fa_7_105_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$273 final_adder.U$$272/A final_adder.U$$161/X final_adder.U$$163/X
+ VGND VGND VPWR VPWR final_adder.U$$273/X sky130_fd_sc_hd__a21o_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$112 U$$934/A1 U$$4/X U$$799/A1 U$$5/X VGND VGND VPWR VPWR U$$113/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$284 final_adder.U$$284/A final_adder.U$$284/B VGND VGND VPWR VPWR
+ final_adder.U$$334/B sky130_fd_sc_hd__and2_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$123 U$$123/A _617_/Q VGND VGND VPWR VPWR U$$123/X sky130_fd_sc_hd__xor2_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$295 final_adder.U$$294/A final_adder.U$$205/X final_adder.U$$207/X
+ VGND VGND VPWR VPWR final_adder.U$$295/X sky130_fd_sc_hd__a21o_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$134 U$$819/A1 U$$4/X U$$134/B1 U$$5/X VGND VGND VPWR VPWR U$$135/A sky130_fd_sc_hd__a22o_1
XFILLER_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$145 U$$8/A1 U$$141/X U$$8/B1 U$$142/X VGND VGND VPWR VPWR U$$146/A sky130_fd_sc_hd__a22o_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_533_ _535_/CLK _533_/D VGND VGND VPWR VPWR _533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_3 dadda_fa_3_25_3/A dadda_fa_3_25_3/B dadda_fa_3_25_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_26_1/B dadda_fa_4_25_2/CIN sky130_fd_sc_hd__fa_2
XU$$156 U$$156/A U$$274/A VGND VGND VPWR VPWR U$$156/X sky130_fd_sc_hd__xor2_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$167 U$$28/B1 U$$141/X U$$32/A1 U$$142/X VGND VGND VPWR VPWR U$$168/A sky130_fd_sc_hd__a22o_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$178 U$$178/A U$$262/B VGND VGND VPWR VPWR U$$178/X sky130_fd_sc_hd__xor2_1
XFILLER_72_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$189 U$$52/A1 U$$141/X U$$54/A1 U$$142/X VGND VGND VPWR VPWR U$$190/A sky130_fd_sc_hd__a22o_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ _464_/CLK _464_/D VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_395_ _537_/CLK _395_/D VGND VGND VPWR VPWR _395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_92_0 dadda_fa_6_92_0/A dadda_fa_6_92_0/B dadda_fa_6_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_93_0/B dadda_fa_7_92_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$690 U$$688/B _625_/Q _626_/Q U$$685/Y VGND VGND VPWR VPWR U$$690/X sky130_fd_sc_hd__a22o_4
XFILLER_182_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_80_8 U$$4290/X U$$4423/X VGND VGND VPWR VPWR dadda_fa_2_81_3/B dadda_fa_3_80_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_118_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_72_5 U$$4008/X U$$4141/X U$$4274/X VGND VGND VPWR VPWR dadda_fa_2_73_2/A
+ dadda_fa_2_72_5/A sky130_fd_sc_hd__fa_2
XFILLER_150_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_65_4 U$$4127/X U$$4260/X U$$4393/X VGND VGND VPWR VPWR dadda_fa_2_66_1/CIN
+ dadda_fa_2_65_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_140_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_58_3 U$$2783/X U$$2916/X U$$3049/X VGND VGND VPWR VPWR dadda_fa_2_59_1/B
+ dadda_fa_2_58_4/B sky130_fd_sc_hd__fa_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_35_2 dadda_fa_4_35_2/A dadda_fa_4_35_2/B dadda_fa_4_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/CIN dadda_fa_5_35_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_1 dadda_fa_4_28_1/A dadda_fa_4_28_1/B dadda_fa_4_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/B dadda_fa_5_28_1/B sky130_fd_sc_hd__fa_2
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_180_ _336_/CLK _180_/D VGND VGND VPWR VPWR _180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4405 U$$4405/A U$$4405/B VGND VGND VPWR VPWR U$$4405/X sky130_fd_sc_hd__xor2_4
XU$$4416 _564_/Q U$$4388/X _565_/Q U$$4389/X VGND VGND VPWR VPWR U$$4417/A sky130_fd_sc_hd__a22o_2
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_60_3 U$$1324/X U$$1457/X U$$1590/X VGND VGND VPWR VPWR dadda_fa_1_61_7/A
+ dadda_fa_1_60_8/CIN sky130_fd_sc_hd__fa_2
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4427 U$$4427/A U$$4427/B VGND VGND VPWR VPWR U$$4427/X sky130_fd_sc_hd__xor2_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4438 U$$4438/A1 U$$4388/X _576_/Q U$$4389/X VGND VGND VPWR VPWR U$$4439/A sky130_fd_sc_hd__a22o_1
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4449 U$$4449/A U$$4449/B VGND VGND VPWR VPWR U$$4449/X sky130_fd_sc_hd__xor2_2
Xdadda_ha_3_17_1 U$$440/X U$$573/X VGND VGND VPWR VPWR dadda_fa_4_18_1/CIN dadda_ha_3_17_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3704 U$$3702/B U$$3699/A _670_/Q U$$3699/Y VGND VGND VPWR VPWR U$$3704/X sky130_fd_sc_hd__a22o_4
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3715 _556_/Q U$$3783/A2 U$$975/B1 U$$3783/B2 VGND VGND VPWR VPWR U$$3716/A sky130_fd_sc_hd__a22o_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3726 U$$3726/A U$$3784/B VGND VGND VPWR VPWR U$$3726/X sky130_fd_sc_hd__xor2_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3737 U$$4285/A1 U$$3795/A2 U$$4424/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3738/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_1 input180/X dadda_fa_3_30_1/B dadda_fa_3_30_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_31_0/CIN dadda_fa_4_30_2/A sky130_fd_sc_hd__fa_1
XU$$3748 U$$3748/A U$$3784/B VGND VGND VPWR VPWR U$$3748/X sky130_fd_sc_hd__xor2_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3759 _578_/Q U$$3783/A2 U$$4446/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3760/A sky130_fd_sc_hd__a22o_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_0 U$$319/X U$$452/X U$$585/X VGND VGND VPWR VPWR dadda_fa_4_24_0/B
+ dadda_fa_4_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_72_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_516_ _518_/CLK _516_/D VGND VGND VPWR VPWR _516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ _447_/CLK _447_/D VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_378_ _509_/CLK _378_/D VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_82_4 dadda_fa_2_82_4/A dadda_fa_2_82_4/B dadda_fa_2_82_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/CIN dadda_fa_3_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_75_3 dadda_fa_2_75_3/A dadda_fa_2_75_3/B dadda_fa_2_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/B dadda_fa_3_75_3/B sky130_fd_sc_hd__fa_2
XFILLER_123_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_2 dadda_fa_2_68_2/A dadda_fa_2_68_2/B dadda_fa_2_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/A dadda_fa_3_68_3/A sky130_fd_sc_hd__fa_2
XFILLER_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_45_1 dadda_fa_5_45_1/A dadda_fa_5_45_1/B dadda_fa_5_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/B dadda_fa_7_45_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_38_0 dadda_fa_5_38_0/A dadda_fa_5_38_0/B dadda_fa_5_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/A dadda_fa_6_38_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_112_0 dadda_fa_5_112_0/A dadda_fa_5_112_0/B dadda_fa_5_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/A dadda_fa_6_112_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_70_2 U$$3073/X U$$3206/X U$$3339/X VGND VGND VPWR VPWR dadda_fa_2_71_1/A
+ dadda_fa_2_70_4/A sky130_fd_sc_hd__fa_2
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_63_1 U$$2793/X U$$2926/X U$$3059/X VGND VGND VPWR VPWR dadda_fa_2_64_0/CIN
+ dadda_fa_2_63_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_8_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_40_0 dadda_fa_4_40_0/A dadda_fa_4_40_0/B dadda_fa_4_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/A dadda_fa_5_40_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_0 U$$1183/X U$$1316/X U$$1449/X VGND VGND VPWR VPWR dadda_fa_2_57_0/B
+ dadda_fa_2_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1609 U$$4486/A1 U$$1641/A2 U$$787/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1610/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_301_ _303_/CLK _301_/D VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_232_ _499_/CLK hold2/X VGND VGND VPWR VPWR _232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_92_3 dadda_fa_3_92_3/A dadda_fa_3_92_3/B dadda_fa_3_92_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/B dadda_fa_4_92_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_85_2 dadda_fa_3_85_2/A dadda_fa_3_85_2/B dadda_fa_3_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/A dadda_fa_4_85_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_78_1 dadda_fa_3_78_1/A dadda_fa_3_78_1/B dadda_fa_3_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/CIN dadda_fa_4_78_2/A sky130_fd_sc_hd__fa_1
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_55_0 dadda_fa_6_55_0/A dadda_fa_6_55_0/B dadda_fa_6_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_56_0/B dadda_fa_7_55_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater509 U$$1466/B2 VGND VGND VPWR VPWR U$$1474/B2 sky130_fd_sc_hd__buf_12
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4202 U$$4476/A1 U$$4114/X U$$94/A1 U$$4115/X VGND VGND VPWR VPWR U$$4203/A sky130_fd_sc_hd__a22o_1
XU$$4213 U$$4213/A _677_/Q VGND VGND VPWR VPWR U$$4213/X sky130_fd_sc_hd__xor2_1
XFILLER_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4224 _605_/Q U$$4244/A2 U$$4500/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4225/A sky130_fd_sc_hd__a22o_1
XU$$4235 U$$4235/A U$$4246/A VGND VGND VPWR VPWR U$$4235/X sky130_fd_sc_hd__xor2_1
XFILLER_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3501 U$$759/B1 U$$3429/X U$$78/A1 U$$3430/X VGND VGND VPWR VPWR U$$3502/A sky130_fd_sc_hd__a22o_1
XU$$4246 U$$4246/A VGND VGND VPWR VPWR U$$4246/Y sky130_fd_sc_hd__inv_1
XU$$3512 U$$3512/A U$$3536/B VGND VGND VPWR VPWR U$$3512/X sky130_fd_sc_hd__xor2_1
XU$$4257 U$$969/A1 U$$4381/A2 U$$12/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4258/A sky130_fd_sc_hd__a22o_1
XFILLER_133_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3523 _597_/Q U$$3545/A2 _598_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3524/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_114_2 dadda_fa_4_114_2/A dadda_fa_4_114_2/B dadda_ha_3_114_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_115_0/CIN dadda_fa_5_114_1/CIN sky130_fd_sc_hd__fa_1
XU$$4268 U$$4268/A U$$4332/B VGND VGND VPWR VPWR U$$4268/X sky130_fd_sc_hd__xor2_1
XU$$4279 _564_/Q U$$4377/A2 _565_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4280/A sky130_fd_sc_hd__a22o_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3534 U$$3534/A U$$3536/B VGND VGND VPWR VPWR U$$3534/X sky130_fd_sc_hd__xor2_1
XU$$3545 U$$942/A1 U$$3545/A2 U$$4506/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3546/A
+ sky130_fd_sc_hd__a22o_1
XU$$2800 _578_/Q U$$2868/A2 U$$3624/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2801/A sky130_fd_sc_hd__a22o_1
XU$$2811 U$$2811/A U$$2871/B VGND VGND VPWR VPWR U$$2811/X sky130_fd_sc_hd__xor2_2
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3556 U$$3556/A U$$3561/A VGND VGND VPWR VPWR U$$3556/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_107_1 dadda_fa_4_107_1/A dadda_fa_4_107_1/B dadda_fa_4_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/B dadda_fa_5_107_1/B sky130_fd_sc_hd__fa_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2822 _589_/Q U$$2870/A2 _590_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2823/A sky130_fd_sc_hd__a22o_1
XFILLER_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3567 U$$3565/B _667_/Q _668_/Q U$$3562/Y VGND VGND VPWR VPWR U$$3567/X sky130_fd_sc_hd__a22o_4
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2833 U$$2833/A U$$2871/B VGND VGND VPWR VPWR U$$2833/X sky130_fd_sc_hd__xor2_1
XU$$3578 U$$16/A1 U$$3678/A2 U$$975/B1 U$$3678/B2 VGND VGND VPWR VPWR U$$3579/A sky130_fd_sc_hd__a22o_1
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2844 U$$787/B1 U$$2868/A2 _601_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2845/A sky130_fd_sc_hd__a22o_1
XU$$3589 U$$3589/A U$$3625/B VGND VGND VPWR VPWR U$$3589/X sky130_fd_sc_hd__xor2_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2855 U$$2855/A _657_/Q VGND VGND VPWR VPWR U$$2855/X sky130_fd_sc_hd__xor2_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2866 _611_/Q U$$2870/A2 U$$950/A1 U$$2870/B2 VGND VGND VPWR VPWR U$$2867/A sky130_fd_sc_hd__a22o_1
XFILLER_61_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2877 _657_/Q VGND VGND VPWR VPWR U$$2877/Y sky130_fd_sc_hd__inv_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2888 U$$2888/A U$$2996/B VGND VGND VPWR VPWR U$$2888/X sky130_fd_sc_hd__xor2_1
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2899 U$$22/A1 U$$2975/A2 U$$4271/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2900/A sky130_fd_sc_hd__a22o_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_80_1 dadda_fa_2_80_1/A dadda_fa_2_80_1/B dadda_fa_2_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_0/CIN dadda_fa_3_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_73_0 dadda_fa_2_73_0/A dadda_fa_2_73_0/B dadda_fa_2_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/B dadda_fa_3_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_64_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_95_1 dadda_fa_4_95_1/A dadda_fa_4_95_1/B dadda_fa_4_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/B dadda_fa_5_95_1/B sky130_fd_sc_hd__fa_2
XFILLER_180_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_72_0 dadda_fa_7_72_0/A dadda_fa_7_72_0/B dadda_fa_7_72_0/CIN VGND VGND
+ VPWR VPWR _497_/D _368_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_88_0 dadda_fa_4_88_0/A dadda_fa_4_88_0/B dadda_fa_4_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/A dadda_fa_5_88_1/A sky130_fd_sc_hd__fa_1
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_109_3 U$$4348/X U$$4481/X input139/X VGND VGND VPWR VPWR dadda_fa_4_110_1/B
+ dadda_fa_4_109_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput370 _255_/Q VGND VGND VPWR VPWR o[87] sky130_fd_sc_hd__buf_2
XFILLER_156_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput381 _265_/Q VGND VGND VPWR VPWR o[97] sky130_fd_sc_hd__buf_2
XFILLER_156_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2107 U$$2790/B1 U$$2117/A2 U$$876/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2108/A
+ sky130_fd_sc_hd__a22o_1
XU$$2118 U$$2118/A U$$2118/B VGND VGND VPWR VPWR U$$2118/X sky130_fd_sc_hd__xor2_1
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2129 U$$759/A1 U$$2059/X U$$759/B1 U$$2060/X VGND VGND VPWR VPWR U$$2130/A sky130_fd_sc_hd__a22o_1
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1406 U$$4283/A1 U$$1474/A2 U$$38/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1407/A sky130_fd_sc_hd__a22o_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1417 U$$1417/A U$$1461/B VGND VGND VPWR VPWR U$$1417/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1428 U$$58/A1 U$$1472/A2 U$$60/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1429/A sky130_fd_sc_hd__a22o_1
XU$$1439 U$$1439/A U$$1505/B VGND VGND VPWR VPWR U$$1439/X sky130_fd_sc_hd__xor2_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_215_ _480_/CLK _215_/D VGND VGND VPWR VPWR _215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_90_0 dadda_fa_3_90_0/A dadda_fa_3_90_0/B dadda_fa_3_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/B dadda_fa_4_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_52_5 dadda_fa_2_52_5/A dadda_fa_2_52_5/B dadda_fa_2_52_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_2/A dadda_fa_4_52_0/A sky130_fd_sc_hd__fa_2
XFILLER_39_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4010 U$$4010/A U$$4044/B VGND VGND VPWR VPWR U$$4010/X sky130_fd_sc_hd__xor2_1
XFILLER_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4021 U$$4156/B1 U$$4045/A2 _573_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$4022/A sky130_fd_sc_hd__a22o_1
XU$$4032 U$$4032/A U$$4044/B VGND VGND VPWR VPWR U$$4032/X sky130_fd_sc_hd__xor2_1
XU$$4043 U$$70/A1 U$$4045/A2 U$$72/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$4044/A sky130_fd_sc_hd__a22o_1
XU$$4054 U$$4054/A U$$4058/B VGND VGND VPWR VPWR U$$4054/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_4 dadda_fa_2_45_4/A dadda_fa_2_45_4/B dadda_fa_2_45_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/CIN dadda_fa_3_45_3/CIN sky130_fd_sc_hd__fa_1
XU$$3320 _564_/Q U$$3396/A2 _565_/Q U$$3396/B2 VGND VGND VPWR VPWR U$$3321/A sky130_fd_sc_hd__a22o_1
XFILLER_47_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4065 U$$4476/A1 U$$4107/A2 U$$94/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4066/A sky130_fd_sc_hd__a22o_1
XU$$4076 U$$4076/A U$$4109/A VGND VGND VPWR VPWR U$$4076/X sky130_fd_sc_hd__xor2_1
XU$$3331 U$$3331/A U$$3413/B VGND VGND VPWR VPWR U$$3331/X sky130_fd_sc_hd__xor2_1
XU$$3342 U$$4438/A1 U$$3396/A2 U$$4303/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3343/A
+ sky130_fd_sc_hd__a22o_1
XU$$4087 _605_/Q U$$4107/A2 U$$4500/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4088/A sky130_fd_sc_hd__a22o_1
XU$$3353 U$$3353/A U$$3403/B VGND VGND VPWR VPWR U$$3353/X sky130_fd_sc_hd__xor2_1
XU$$4098 U$$4098/A U$$4109/A VGND VGND VPWR VPWR U$$4098/X sky130_fd_sc_hd__xor2_1
XU$$3364 _586_/Q U$$3292/X _587_/Q U$$3293/X VGND VGND VPWR VPWR U$$3365/A sky130_fd_sc_hd__a22o_1
XFILLER_19_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_38_3 U$$2344/X U$$2477/X U$$2610/X VGND VGND VPWR VPWR dadda_fa_3_39_1/B
+ dadda_fa_3_38_3/B sky130_fd_sc_hd__fa_1
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2630 U$$2630/A U$$2710/B VGND VGND VPWR VPWR U$$2630/X sky130_fd_sc_hd__xor2_1
XU$$3375 U$$3375/A U$$3413/B VGND VGND VPWR VPWR U$$3375/X sky130_fd_sc_hd__xor2_1
XFILLER_179_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2641 U$$4285/A1 U$$2667/A2 U$$3191/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2642/A
+ sky130_fd_sc_hd__a22o_1
XU$$3386 U$$98/A1 U$$3412/A2 U$$98/B1 U$$3412/B2 VGND VGND VPWR VPWR U$$3387/A sky130_fd_sc_hd__a22o_1
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2652 U$$2652/A U$$2698/B VGND VGND VPWR VPWR U$$2652/X sky130_fd_sc_hd__xor2_1
XU$$3397 U$$3397/A U$$3397/B VGND VGND VPWR VPWR U$$3397/X sky130_fd_sc_hd__xor2_1
XU$$2663 _578_/Q U$$2729/A2 U$$4446/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2664/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2674 U$$2674/A U$$2698/B VGND VGND VPWR VPWR U$$2674/X sky130_fd_sc_hd__xor2_1
XU$$1940 U$$979/B1 U$$2036/A2 U$$4271/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1941/A
+ sky130_fd_sc_hd__a22o_1
XU$$2685 U$$902/B1 U$$2729/A2 U$$84/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2686/A sky130_fd_sc_hd__a22o_1
XU$$1951 U$$1951/A U$$1991/B VGND VGND VPWR VPWR U$$1951/X sky130_fd_sc_hd__xor2_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2696 U$$2696/A U$$2698/B VGND VGND VPWR VPWR U$$2696/X sky130_fd_sc_hd__xor2_1
XU$$1962 U$$4291/A1 U$$1922/X U$$868/A1 U$$1923/X VGND VGND VPWR VPWR U$$1963/A sky130_fd_sc_hd__a22o_1
XFILLER_178_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1973 U$$1973/A U$$1991/B VGND VGND VPWR VPWR U$$1973/X sky130_fd_sc_hd__xor2_1
XU$$1984 U$$3489/B1 U$$2036/A2 U$$3217/B1 U$$2036/B2 VGND VGND VPWR VPWR U$$1985/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1995 U$$1995/A U$$2021/B VGND VGND VPWR VPWR U$$1995/X sky130_fd_sc_hd__xor2_1
XFILLER_193_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_732__784 VGND VGND VPWR VPWR _732__784/HI U$$2335/A1 sky130_fd_sc_hd__conb_1
XFILLER_131_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput109 b[4] VGND VGND VPWR VPWR _556_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$603 final_adder.U$$730/A final_adder.U$$730/B final_adder.U$$603/B1
+ VGND VGND VPWR VPWR final_adder.U$$731/B sky130_fd_sc_hd__a21o_1
XFILLER_5_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$625 final_adder.U$$625/A final_adder.U$$625/B VGND VGND VPWR VPWR
+ _171_/D sky130_fd_sc_hd__xor2_4
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$636 final_adder.U$$636/A final_adder.U$$636/B VGND VGND VPWR VPWR
+ hold4/A sky130_fd_sc_hd__xor2_1
XFILLER_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$647 final_adder.U$$647/A final_adder.U$$647/B VGND VGND VPWR VPWR
+ _193_/D sky130_fd_sc_hd__xor2_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$658 final_adder.U$$658/A final_adder.U$$658/B VGND VGND VPWR VPWR
+ _204_/D sky130_fd_sc_hd__xor2_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$669 final_adder.U$$669/A final_adder.U$$669/B VGND VGND VPWR VPWR
+ _215_/D sky130_fd_sc_hd__xor2_1
XU$$508 U$$508/A U$$547/A VGND VGND VPWR VPWR U$$508/X sky130_fd_sc_hd__xor2_1
XU$$519 U$$928/B1 U$$545/A2 _603_/Q U$$416/X VGND VGND VPWR VPWR U$$520/A sky130_fd_sc_hd__a22o_1
XFILLER_38_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$80 U$$80/A1 U$$4/X U$$82/A1 U$$5/X VGND VGND VPWR VPWR U$$81/A sky130_fd_sc_hd__a22o_1
XFILLER_53_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$91 U$$91/A U$$3/A VGND VGND VPWR VPWR U$$91/X sky130_fd_sc_hd__xor2_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_0 U$$3413/X U$$3546/X U$$3679/X VGND VGND VPWR VPWR dadda_fa_4_108_0/B
+ dadda_fa_4_107_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_55_3 dadda_fa_3_55_3/A dadda_fa_3_55_3/B dadda_fa_3_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/B dadda_fa_4_55_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_681__901 VGND VGND VPWR VPWR _681__901/HI _681__901/LO sky130_fd_sc_hd__conb_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_48_2 dadda_fa_3_48_2/A dadda_fa_3_48_2/B dadda_fa_3_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/A dadda_fa_4_48_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_18_0 dadda_fa_6_18_0/A dadda_fa_6_18_0/B dadda_fa_6_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_19_0/B dadda_fa_7_18_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1203 U$$1203/A _633_/Q VGND VGND VPWR VPWR U$$1203/X sky130_fd_sc_hd__xor2_1
XU$$1214 U$$940/A1 U$$1100/X U$$942/A1 U$$1101/X VGND VGND VPWR VPWR U$$1215/A sky130_fd_sc_hd__a22o_1
XU$$1225 U$$1225/A _633_/Q VGND VGND VPWR VPWR U$$1225/X sky130_fd_sc_hd__xor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1236 _635_/Q U$$1236/B VGND VGND VPWR VPWR U$$1236/X sky130_fd_sc_hd__and2_1
XU$$1247 U$$12/B1 U$$1237/X U$$14/B1 U$$1238/X VGND VGND VPWR VPWR U$$1248/A sky130_fd_sc_hd__a22o_1
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1258 U$$1258/A U$$1336/B VGND VGND VPWR VPWR U$$1258/X sky130_fd_sc_hd__xor2_1
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1269 U$$4283/A1 U$$1341/A2 U$$38/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1270/A sky130_fd_sc_hd__a22o_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_716__768 VGND VGND VPWR VPWR _716__768/HI U$$1367/B1 sky130_fd_sc_hd__conb_1
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_50_2 dadda_fa_2_50_2/A dadda_fa_2_50_2/B dadda_fa_2_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/A dadda_fa_3_50_3/A sky130_fd_sc_hd__fa_2
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_43_1 U$$2354/X U$$2487/X U$$2620/X VGND VGND VPWR VPWR dadda_fa_3_44_0/CIN
+ dadda_fa_3_43_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_20_0 dadda_fa_5_20_0/A dadda_fa_5_20_0/B dadda_fa_5_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/A dadda_fa_6_20_0/CIN sky130_fd_sc_hd__fa_1
XU$$3150 _661_/Q VGND VGND VPWR VPWR U$$3150/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_0 U$$744/X U$$877/X U$$1010/X VGND VGND VPWR VPWR dadda_fa_3_37_0/B
+ dadda_fa_3_36_2/B sky130_fd_sc_hd__fa_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3161 U$$969/A1 U$$3241/A2 U$$12/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3162/A sky130_fd_sc_hd__a22o_1
XU$$3172 U$$3172/A U$$3244/B VGND VGND VPWR VPWR U$$3172/X sky130_fd_sc_hd__xor2_1
XU$$3183 _564_/Q U$$3243/A2 _565_/Q U$$3243/B2 VGND VGND VPWR VPWR U$$3184/A sky130_fd_sc_hd__a22o_1
XU$$3194 U$$3194/A U$$3224/B VGND VGND VPWR VPWR U$$3194/X sky130_fd_sc_hd__xor2_1
XFILLER_179_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2460 U$$2460/A _651_/Q VGND VGND VPWR VPWR U$$2460/X sky130_fd_sc_hd__xor2_1
XU$$2471 U$$2469/B _651_/Q _652_/Q U$$2466/Y VGND VGND VPWR VPWR U$$2471/X sky130_fd_sc_hd__a22o_4
XU$$2482 U$$16/A1 U$$2574/A2 U$$18/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2483/A sky130_fd_sc_hd__a22o_1
XU$$2493 U$$2493/A U$$2533/B VGND VGND VPWR VPWR U$$2493/X sky130_fd_sc_hd__xor2_1
XFILLER_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1770 _611_/Q U$$1770/A2 _612_/Q U$$1770/B2 VGND VGND VPWR VPWR U$$1771/A sky130_fd_sc_hd__a22o_1
XFILLER_50_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1781 U$$1781/A VGND VGND VPWR VPWR U$$1781/Y sky130_fd_sc_hd__inv_1
XFILLER_148_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1792 U$$1792/A U$$1918/A VGND VGND VPWR VPWR U$$1792/X sky130_fd_sc_hd__xor2_1
XFILLER_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput80 b[23] VGND VGND VPWR VPWR _575_/D sky130_fd_sc_hd__buf_2
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput91 b[33] VGND VGND VPWR VPWR _585_/D sky130_fd_sc_hd__buf_2
XFILLER_66_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_88_3 U$$2843/X U$$2976/X U$$3109/X VGND VGND VPWR VPWR dadda_fa_2_89_4/B
+ dadda_fa_2_88_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_65_2 dadda_fa_4_65_2/A dadda_fa_4_65_2/B dadda_fa_4_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/CIN dadda_fa_5_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_58_1 dadda_fa_4_58_1/A dadda_fa_4_58_1/B dadda_fa_4_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/B dadda_fa_5_58_1/B sky130_fd_sc_hd__fa_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$411 final_adder.U$$328/B final_adder.U$$654/B final_adder.U$$273/X
+ VGND VGND VPWR VPWR final_adder.U$$658/B sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_35_0 dadda_fa_7_35_0/A dadda_fa_7_35_0/B dadda_fa_7_35_0/CIN VGND VGND
+ VPWR VPWR _460_/D _331_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$433 final_adder.U$$316/X final_adder.U$$742/B final_adder.U$$317/X
+ VGND VGND VPWR VPWR final_adder.U$$746/B sky130_fd_sc_hd__a21o_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$455 final_adder.U$$278/B final_adder.U$$666/B final_adder.U$$173/X
+ VGND VGND VPWR VPWR final_adder.U$$668/B sky130_fd_sc_hd__a21o_1
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$305 U$$305/A U$$391/B VGND VGND VPWR VPWR U$$305/X sky130_fd_sc_hd__xor2_1
X_706__926 VGND VGND VPWR VPWR _706__926/HI _706__926/LO sky130_fd_sc_hd__conb_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater670 U$$630/A1 VGND VGND VPWR VPWR U$$82/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$477 final_adder.U$$300/B final_adder.U$$710/B final_adder.U$$217/X
+ VGND VGND VPWR VPWR final_adder.U$$712/B sky130_fd_sc_hd__a21o_1
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$316 _569_/Q U$$278/X _570_/Q U$$279/X VGND VGND VPWR VPWR U$$317/A sky130_fd_sc_hd__a22o_1
Xrepeater681 U$$4045/B1 VGND VGND VPWR VPWR U$$759/A1 sky130_fd_sc_hd__buf_12
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$327 U$$327/A U$$357/B VGND VGND VPWR VPWR U$$327/X sky130_fd_sc_hd__xor2_1
Xrepeater692 _581_/Q VGND VGND VPWR VPWR U$$66/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$499 final_adder.U$$626/A final_adder.U$$626/B final_adder.U$$499/B1
+ VGND VGND VPWR VPWR final_adder.U$$627/B sky130_fd_sc_hd__a21o_1
XU$$338 U$$64/A1 U$$278/X U$$66/A1 U$$279/X VGND VGND VPWR VPWR U$$339/A sky130_fd_sc_hd__a22o_1
XFILLER_123_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$349 U$$349/A U$$391/B VGND VGND VPWR VPWR U$$349/X sky130_fd_sc_hd__xor2_1
X_480_ _480_/CLK _480_/D VGND VGND VPWR VPWR _480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_60_1 dadda_fa_3_60_1/A dadda_fa_3_60_1/B dadda_fa_3_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/CIN dadda_fa_4_60_2/A sky130_fd_sc_hd__fa_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_53_0 dadda_fa_3_53_0/A dadda_fa_3_53_0/B dadda_fa_3_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/B dadda_fa_4_53_1/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_0_69_0 U$$410/Y U$$544/X U$$677/X VGND VGND VPWR VPWR dadda_fa_1_70_6/A
+ dadda_fa_1_69_7/CIN sky130_fd_sc_hd__fa_2
XFILLER_48_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$850 U$$987/A1 U$$928/A2 U$$28/B1 U$$928/B2 VGND VGND VPWR VPWR U$$851/A sky130_fd_sc_hd__a22o_1
X_678_ _678_/CLK _678_/D VGND VGND VPWR VPWR _678_/Q sky130_fd_sc_hd__dfxtp_1
XU$$861 U$$861/A U$$959/A VGND VGND VPWR VPWR U$$861/X sky130_fd_sc_hd__xor2_1
XU$$1000 U$$999/X U$$992/B VGND VGND VPWR VPWR U$$1000/X sky130_fd_sc_hd__xor2_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$872 U$$50/A1 U$$910/A2 U$$50/B1 U$$910/B2 VGND VGND VPWR VPWR U$$873/A sky130_fd_sc_hd__a22o_1
XU$$1011 U$$2790/B1 U$$999/A2 U$$876/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1012/A sky130_fd_sc_hd__a22o_1
XU$$1022 U$$1022/A U$$992/B VGND VGND VPWR VPWR U$$1022/X sky130_fd_sc_hd__xor2_1
XU$$883 U$$883/A U$$903/B VGND VGND VPWR VPWR U$$883/X sky130_fd_sc_hd__xor2_1
XFILLER_32_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1033 U$$74/A1 U$$1093/A2 U$$76/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1034/A sky130_fd_sc_hd__a22o_1
XU$$894 U$$72/A1 U$$910/A2 U$$74/A1 U$$910/B2 VGND VGND VPWR VPWR U$$895/A sky130_fd_sc_hd__a22o_1
XU$$1044 U$$1044/A U$$992/B VGND VGND VPWR VPWR U$$1044/X sky130_fd_sc_hd__xor2_1
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1055 U$$94/B1 U$$1093/A2 U$$98/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1056/A sky130_fd_sc_hd__a22o_1
XFILLER_16_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1066 U$$1066/A U$$998/B VGND VGND VPWR VPWR U$$1066/X sky130_fd_sc_hd__xor2_1
XU$$1077 U$$940/A1 U$$963/X U$$942/A1 U$$964/X VGND VGND VPWR VPWR U$$1078/A sky130_fd_sc_hd__a22o_1
XFILLER_149_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1088 U$$1088/A _631_/Q VGND VGND VPWR VPWR U$$1088/X sky130_fd_sc_hd__xor2_1
XFILLER_188_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1099 _633_/Q U$$1099/B VGND VGND VPWR VPWR U$$1099/X sky130_fd_sc_hd__and2_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_110_0 dadda_fa_7_110_0/A dadda_fa_7_110_0/B dadda_fa_7_110_0/CIN VGND
+ VGND VPWR VPWR _535_/D _406_/D sky130_fd_sc_hd__fa_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_98_2 U$$3129/X U$$3262/X U$$3395/X VGND VGND VPWR VPWR dadda_fa_3_99_1/B
+ dadda_fa_3_98_3/A sky130_fd_sc_hd__fa_1
XFILLER_176_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_75_1 dadda_fa_5_75_1/A dadda_fa_5_75_1/B dadda_fa_5_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/B dadda_fa_7_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_68_0 dadda_fa_5_68_0/A dadda_fa_5_68_0/B dadda_fa_5_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/A dadda_fa_6_68_0/CIN sky130_fd_sc_hd__fa_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_8 dadda_fa_1_67_8/A dadda_fa_1_67_8/B dadda_fa_1_67_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_3/A dadda_fa_3_67_0/A sky130_fd_sc_hd__fa_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_844__896 VGND VGND VPWR VPWR _844__896/HI U$$828/A1 sky130_fd_sc_hd__conb_1
XFILLER_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_7_0 dadda_fa_6_7_0/A dadda_fa_6_7_0/B dadda_fa_6_7_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_8_0/B dadda_fa_7_7_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2290 _597_/Q U$$2326/A2 _598_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2291/A sky130_fd_sc_hd__a22o_1
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_738__790 VGND VGND VPWR VPWR _738__790/HI U$$2737/B1 sky130_fd_sc_hd__conb_1
XFILLER_191_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_93_1 U$$2454/X U$$2587/X U$$2720/X VGND VGND VPWR VPWR dadda_fa_2_94_5/B
+ dadda_fa_3_93_0/A sky130_fd_sc_hd__fa_2
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_70_0 dadda_fa_4_70_0/A dadda_fa_4_70_0/B dadda_fa_4_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/A dadda_fa_5_70_1/A sky130_fd_sc_hd__fa_1
XFILLER_2_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_86_0 _688__908/HI U$$1642/X U$$1775/X VGND VGND VPWR VPWR dadda_fa_2_87_2/CIN
+ dadda_fa_2_86_4/B sky130_fd_sc_hd__fa_2
XFILLER_150_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_106_1 U$$3278/X U$$3411/X VGND VGND VPWR VPWR dadda_fa_3_107_3/CIN dadda_fa_4_106_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$230 final_adder.U$$725/A final_adder.U$$724/A VGND VGND VPWR VPWR
+ final_adder.U$$306/A sky130_fd_sc_hd__and2_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3908 _584_/Q U$$3840/X _585_/Q U$$3841/X VGND VGND VPWR VPWR U$$3909/A sky130_fd_sc_hd__a22o_1
XFILLER_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$241 final_adder.U$$735/A final_adder.U$$607/B1 final_adder.U$$241/B1
+ VGND VGND VPWR VPWR final_adder.U$$241/X sky130_fd_sc_hd__a21o_1
X_601_ _601_/CLK _601_/D VGND VGND VPWR VPWR _601_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3919 U$$3919/A U$$3969/B VGND VGND VPWR VPWR U$$3919/X sky130_fd_sc_hd__xor2_1
XFILLER_58_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$252 final_adder.U$$747/A final_adder.U$$746/A VGND VGND VPWR VPWR
+ final_adder.U$$252/X sky130_fd_sc_hd__and2_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$263 final_adder.U$$262/A final_adder.U$$141/X final_adder.U$$143/X
+ VGND VGND VPWR VPWR final_adder.U$$263/X sky130_fd_sc_hd__a21o_1
XU$$102 U$$924/A1 U$$4/X U$$926/A1 U$$5/X VGND VGND VPWR VPWR U$$103/A sky130_fd_sc_hd__a22o_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$274 final_adder.U$$274/A final_adder.U$$274/B VGND VGND VPWR VPWR
+ final_adder.U$$328/A sky130_fd_sc_hd__and2_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$113 U$$113/A _617_/Q VGND VGND VPWR VPWR U$$113/X sky130_fd_sc_hd__xor2_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$285 final_adder.U$$284/A final_adder.U$$185/X final_adder.U$$187/X
+ VGND VGND VPWR VPWR final_adder.U$$285/X sky130_fd_sc_hd__a21o_1
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$124 U$$946/A1 U$$4/X U$$948/A1 U$$5/X VGND VGND VPWR VPWR U$$125/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$296 final_adder.U$$296/A final_adder.U$$296/B VGND VGND VPWR VPWR
+ final_adder.U$$340/B sky130_fd_sc_hd__and2_1
X_532_ _532_/CLK _532_/D VGND VGND VPWR VPWR _532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$135 U$$135/A U$$89/B VGND VGND VPWR VPWR U$$135/X sky130_fd_sc_hd__xor2_1
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$146 U$$146/A U$$242/B VGND VGND VPWR VPWR U$$146/X sky130_fd_sc_hd__xor2_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$157 U$$842/A1 U$$141/X U$$22/A1 U$$142/X VGND VGND VPWR VPWR U$$158/A sky130_fd_sc_hd__a22o_1
XFILLER_45_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$168 U$$168/A U$$262/B VGND VGND VPWR VPWR U$$168/X sky130_fd_sc_hd__xor2_1
XFILLER_45_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$179 _569_/Q U$$141/X _570_/Q U$$142/X VGND VGND VPWR VPWR U$$180/A sky130_fd_sc_hd__a22o_1
X_463_ _463_/CLK _463_/D VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_394_ _535_/CLK _394_/D VGND VGND VPWR VPWR _394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_85_0 dadda_fa_6_85_0/A dadda_fa_6_85_0/B dadda_fa_6_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_86_0/B dadda_fa_7_85_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_787__839 VGND VGND VPWR VPWR _787__839/HI U$$4419/B sky130_fd_sc_hd__conb_1
XFILLER_49_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$680 U$$952/B1 U$$682/A2 U$$956/A1 U$$553/X VGND VGND VPWR VPWR U$$681/A sky130_fd_sc_hd__a22o_1
XU$$691 U$$691/A1 U$$817/A2 _552_/Q U$$785/B2 VGND VGND VPWR VPWR U$$692/A sky130_fd_sc_hd__a22o_2
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_72_6 U$$4407/X input226/X dadda_fa_1_72_6/CIN VGND VGND VPWR VPWR dadda_fa_2_73_2/B
+ dadda_fa_2_72_5/B sky130_fd_sc_hd__fa_2
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_65_5 input218/X dadda_fa_1_65_5/B dadda_fa_1_65_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_66_2/A dadda_fa_2_65_5/A sky130_fd_sc_hd__fa_1
XFILLER_58_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_58_4 U$$3182/X U$$3315/X U$$3448/X VGND VGND VPWR VPWR dadda_fa_2_59_1/CIN
+ dadda_fa_2_58_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk _632_/CLK VGND VGND VPWR VPWR _621_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_28_2 dadda_fa_4_28_2/A dadda_fa_4_28_2/B dadda_fa_4_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/CIN dadda_fa_5_28_1/CIN sky130_fd_sc_hd__fa_2
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4406 _559_/Q U$$4388/X _560_/Q U$$4389/X VGND VGND VPWR VPWR U$$4407/A sky130_fd_sc_hd__a22o_1
XFILLER_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4417 U$$4417/A U$$4417/B VGND VGND VPWR VPWR U$$4417/X sky130_fd_sc_hd__xor2_4
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4428 _570_/Q U$$4388/X _571_/Q U$$4389/X VGND VGND VPWR VPWR U$$4429/A sky130_fd_sc_hd__a22o_1
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4439 U$$4439/A U$$4439/B VGND VGND VPWR VPWR U$$4439/X sky130_fd_sc_hd__xor2_1
XFILLER_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3705 U$$3705/A1 U$$3795/A2 U$$4255/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3706/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3716 U$$3716/A U$$3756/B VGND VGND VPWR VPWR U$$3716/X sky130_fd_sc_hd__xor2_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3727 _562_/Q U$$3783/A2 _563_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3728/A sky130_fd_sc_hd__a22o_1
XFILLER_79_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3738 U$$3738/A U$$3756/B VGND VGND VPWR VPWR U$$3738/X sky130_fd_sc_hd__xor2_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3749 U$$735/A1 U$$3783/A2 _574_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3750/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_84_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _644_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_2 dadda_fa_3_30_2/A dadda_fa_3_30_2/B dadda_fa_3_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/A dadda_fa_4_30_2/B sky130_fd_sc_hd__fa_1
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_515_ _515_/CLK _515_/D VGND VGND VPWR VPWR _515_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_3_23_1 U$$718/X U$$851/X U$$984/X VGND VGND VPWR VPWR dadda_fa_4_24_0/CIN
+ dadda_fa_4_23_2/A sky130_fd_sc_hd__fa_2
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_16_0 U$$39/X U$$172/X U$$305/X VGND VGND VPWR VPWR dadda_fa_4_17_1/CIN
+ dadda_fa_4_16_2/B sky130_fd_sc_hd__fa_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_446_ _455_/CLK _446_/D VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_377_ _510_/CLK _377_/D VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_82_5 dadda_fa_2_82_5/A dadda_fa_2_82_5/B dadda_fa_2_82_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_2/A dadda_fa_4_82_0/A sky130_fd_sc_hd__fa_1
XFILLER_79_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_75_4 dadda_fa_2_75_4/A dadda_fa_2_75_4/B dadda_fa_2_75_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/CIN dadda_fa_3_75_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_3 dadda_fa_2_68_3/A dadda_fa_2_68_3/B dadda_fa_2_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/B dadda_fa_3_68_3/B sky130_fd_sc_hd__fa_1
XFILLER_84_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_38_1 dadda_fa_5_38_1/A dadda_fa_5_38_1/B dadda_fa_5_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/B dadda_fa_7_38_0/A sky130_fd_sc_hd__fa_2
XFILLER_49_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_75_clk _560_/CLK VGND VGND VPWR VPWR _667_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_112_1 dadda_fa_5_112_1/A dadda_fa_5_112_1/B dadda_fa_5_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/B dadda_fa_7_112_0/A sky130_fd_sc_hd__fa_1
XFILLER_146_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_105_0 dadda_fa_5_105_0/A dadda_fa_5_105_0/B dadda_fa_5_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/A dadda_fa_6_105_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_70_3 U$$3472/X U$$3605/X U$$3738/X VGND VGND VPWR VPWR dadda_fa_2_71_1/B
+ dadda_fa_2_70_4/B sky130_fd_sc_hd__fa_1
XFILLER_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_63_2 U$$3192/X U$$3325/X U$$3458/X VGND VGND VPWR VPWR dadda_fa_2_64_1/A
+ dadda_fa_2_63_4/A sky130_fd_sc_hd__fa_2
XFILLER_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_40_1 dadda_fa_4_40_1/A dadda_fa_4_40_1/B dadda_fa_4_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/B dadda_fa_5_40_1/B sky130_fd_sc_hd__fa_1
XFILLER_115_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_56_1 U$$1582/X U$$1715/X U$$1848/X VGND VGND VPWR VPWR dadda_fa_2_57_0/CIN
+ dadda_fa_2_56_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_33_0 dadda_fa_4_33_0/A dadda_fa_4_33_0/B dadda_fa_4_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/A dadda_fa_5_33_1/A sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_66_clk _560_/CLK VGND VGND VPWR VPWR _578_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_49_0 U$$105/X U$$238/X U$$371/X VGND VGND VPWR VPWR dadda_fa_2_50_0/CIN
+ dadda_fa_2_49_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_55_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _327_/CLK _300_/D VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_231_ _499_/CLK _231_/D VGND VGND VPWR VPWR _231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_85_3 dadda_fa_3_85_3/A dadda_fa_3_85_3/B dadda_fa_3_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/B dadda_fa_4_85_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_78_2 dadda_fa_3_78_2/A dadda_fa_3_78_2/B dadda_fa_3_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/A dadda_fa_4_78_2/B sky130_fd_sc_hd__fa_2
XFILLER_85_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_48_0 dadda_fa_6_48_0/A dadda_fa_6_48_0/B dadda_fa_6_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_49_0/B dadda_fa_7_48_0/CIN sky130_fd_sc_hd__fa_2
XU$$4203 U$$4203/A _677_/Q VGND VGND VPWR VPWR U$$4203/X sky130_fd_sc_hd__xor2_1
XU$$4214 U$$787/B1 U$$4244/A2 U$$654/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4215/A sky130_fd_sc_hd__a22o_1
XU$$4225 U$$4225/A U$$4246/A VGND VGND VPWR VPWR U$$4225/X sky130_fd_sc_hd__xor2_1
XFILLER_78_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4236 _611_/Q U$$4244/A2 U$$539/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4237/A sky130_fd_sc_hd__a22o_1
XFILLER_93_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3502 U$$3502/A U$$3561/A VGND VGND VPWR VPWR U$$3502/X sky130_fd_sc_hd__xor2_1
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4247 U$$4247/A VGND VGND VPWR VPWR U$$4247/Y sky130_fd_sc_hd__inv_1
XU$$3513 U$$4335/A1 U$$3545/A2 _593_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3514/A sky130_fd_sc_hd__a22o_1
XU$$4258 U$$4258/A U$$4384/A VGND VGND VPWR VPWR U$$4258/X sky130_fd_sc_hd__xor2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3524 U$$3524/A U$$3536/B VGND VGND VPWR VPWR U$$3524/X sky130_fd_sc_hd__xor2_1
XU$$4269 _559_/Q U$$4381/A2 _560_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4270/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_57_clk _536_/CLK VGND VGND VPWR VPWR _595_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3535 U$$4494/A1 U$$3545/A2 _604_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3536/A sky130_fd_sc_hd__a22o_1
XU$$3546 U$$3546/A _667_/Q VGND VGND VPWR VPWR U$$3546/X sky130_fd_sc_hd__xor2_1
XFILLER_92_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2801 U$$2801/A U$$2839/B VGND VGND VPWR VPWR U$$2801/X sky130_fd_sc_hd__xor2_1
XU$$2812 _584_/Q U$$2870/A2 _585_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2813/A sky130_fd_sc_hd__a22o_1
XU$$3557 U$$4379/A1 U$$3429/X U$$819/A1 U$$3430/X VGND VGND VPWR VPWR U$$3558/A sky130_fd_sc_hd__a22o_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2823 U$$2823/A U$$2871/B VGND VGND VPWR VPWR U$$2823/X sky130_fd_sc_hd__xor2_1
XFILLER_19_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3568 U$$3568/A1 U$$3678/A2 U$$4255/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3569/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_107_2 dadda_fa_4_107_2/A dadda_fa_4_107_2/B dadda_fa_4_107_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/CIN dadda_fa_5_107_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2834 _595_/Q U$$2870/A2 _596_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2835/A sky130_fd_sc_hd__a22o_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3579 U$$3579/A U$$3698/A VGND VGND VPWR VPWR U$$3579/X sky130_fd_sc_hd__xor2_1
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2845 U$$2845/A U$$2871/B VGND VGND VPWR VPWR U$$2845/X sky130_fd_sc_hd__xor2_1
XU$$2856 _606_/Q U$$2870/A2 _607_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2857/A sky130_fd_sc_hd__a22o_1
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2867 U$$2867/A U$$2871/B VGND VGND VPWR VPWR U$$2867/X sky130_fd_sc_hd__xor2_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2878 _658_/Q VGND VGND VPWR VPWR U$$2880/B sky130_fd_sc_hd__inv_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2889 U$$4122/A1 U$$2975/A2 U$$14/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2890/A sky130_fd_sc_hd__a22o_1
XFILLER_18_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _429_/CLK _429_/D VGND VGND VPWR VPWR _429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_80_2 dadda_fa_2_80_2/A dadda_fa_2_80_2/B dadda_fa_2_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/A dadda_fa_3_80_3/A sky130_fd_sc_hd__fa_2
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_73_1 dadda_fa_2_73_1/A dadda_fa_2_73_1/B dadda_fa_2_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/CIN dadda_fa_3_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_50_0 dadda_fa_5_50_0/A dadda_fa_5_50_0/B dadda_fa_5_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/A dadda_fa_6_50_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_66_0 dadda_fa_2_66_0/A dadda_fa_2_66_0/B dadda_fa_2_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/B dadda_fa_3_66_2/B sky130_fd_sc_hd__fa_2
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 a[0] VGND VGND VPWR VPWR _616_/D sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_48_clk _536_/CLK VGND VGND VPWR VPWR _611_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_95_2 dadda_fa_4_95_2/A dadda_fa_4_95_2/B dadda_fa_4_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/CIN dadda_fa_5_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_88_1 dadda_fa_4_88_1/A dadda_fa_4_88_1/B dadda_fa_4_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/B dadda_fa_5_88_1/B sky130_fd_sc_hd__fa_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_65_0 dadda_fa_7_65_0/A dadda_fa_7_65_0/B dadda_fa_7_65_0/CIN VGND VGND
+ VPWR VPWR _490_/D _361_/D sky130_fd_sc_hd__fa_2
XFILLER_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput360 _246_/Q VGND VGND VPWR VPWR o[78] sky130_fd_sc_hd__buf_2
XFILLER_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput371 _256_/Q VGND VGND VPWR VPWR o[88] sky130_fd_sc_hd__buf_2
Xoutput382 _266_/Q VGND VGND VPWR VPWR o[98] sky130_fd_sc_hd__buf_2
XFILLER_120_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _503_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2108 U$$2108/A U$$2118/B VGND VGND VPWR VPWR U$$2108/X sky130_fd_sc_hd__xor2_1
XFILLER_62_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2119 U$$3900/A1 U$$2161/A2 U$$3489/B1 U$$2161/B2 VGND VGND VPWR VPWR U$$2120/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1407 U$$1407/A U$$1461/B VGND VGND VPWR VPWR U$$1407/X sky130_fd_sc_hd__xor2_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1418 U$$48/A1 U$$1472/A2 U$$50/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1419/A sky130_fd_sc_hd__a22o_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1429 U$$1429/A U$$1461/B VGND VGND VPWR VPWR U$$1429/X sky130_fd_sc_hd__xor2_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_214_ _456_/CLK _214_/D VGND VGND VPWR VPWR _214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_90_1 dadda_fa_3_90_1/A dadda_fa_3_90_1/B dadda_fa_3_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/CIN dadda_fa_4_90_2/A sky130_fd_sc_hd__fa_2
XFILLER_100_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_83_0 dadda_fa_3_83_0/A dadda_fa_3_83_0/B dadda_fa_3_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/B dadda_fa_4_83_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_136_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4000 U$$4000/A U$$4058/B VGND VGND VPWR VPWR U$$4000/X sky130_fd_sc_hd__xor2_1
XU$$4011 _567_/Q U$$4107/A2 U$$4424/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4012/A sky130_fd_sc_hd__a22o_1
XFILLER_78_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4022 U$$4022/A U$$4044/B VGND VGND VPWR VPWR U$$4022/X sky130_fd_sc_hd__xor2_1
XU$$4033 U$$4170/A1 U$$4045/A2 U$$4446/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$4034/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4044 U$$4044/A U$$4044/B VGND VGND VPWR VPWR U$$4044/X sky130_fd_sc_hd__xor2_1
XFILLER_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3310 U$$22/A1 U$$3412/A2 _560_/Q U$$3412/B2 VGND VGND VPWR VPWR U$$3311/A sky130_fd_sc_hd__a22o_1
XU$$4055 U$$630/A1 U$$3977/X _590_/Q U$$3978/X VGND VGND VPWR VPWR U$$4056/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_112_0 U$$4354/X U$$4487/X input143/X VGND VGND VPWR VPWR dadda_fa_5_113_0/A
+ dadda_fa_5_112_1/A sky130_fd_sc_hd__fa_2
XU$$4066 U$$4066/A _675_/Q VGND VGND VPWR VPWR U$$4066/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_5 dadda_fa_2_45_5/A dadda_fa_2_45_5/B dadda_fa_2_45_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_2/A dadda_fa_4_45_0/A sky130_fd_sc_hd__fa_2
XU$$3321 U$$3321/A U$$3397/B VGND VGND VPWR VPWR U$$3321/X sky130_fd_sc_hd__xor2_1
XU$$4077 U$$787/B1 U$$4107/A2 U$$654/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4078/A sky130_fd_sc_hd__a22o_1
XU$$3332 U$$4291/A1 U$$3412/A2 U$$46/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3333/A sky130_fd_sc_hd__a22o_1
XU$$3343 U$$3343/A U$$3397/B VGND VGND VPWR VPWR U$$3343/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4088 U$$4088/A U$$4109/A VGND VGND VPWR VPWR U$$4088/X sky130_fd_sc_hd__xor2_1
XU$$3354 _581_/Q U$$3292/X U$$4178/A1 U$$3293/X VGND VGND VPWR VPWR U$$3355/A sky130_fd_sc_hd__a22o_1
XU$$4099 _611_/Q U$$4107/A2 U$$539/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4100/A sky130_fd_sc_hd__a22o_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_38_4 U$$2710/B input188/X dadda_fa_2_38_4/CIN VGND VGND VPWR VPWR dadda_fa_3_39_1/CIN
+ dadda_fa_3_38_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3365 U$$3365/A U$$3403/B VGND VGND VPWR VPWR U$$3365/X sky130_fd_sc_hd__xor2_1
XU$$2620 U$$2620/A U$$2694/B VGND VGND VPWR VPWR U$$2620/X sky130_fd_sc_hd__xor2_1
XFILLER_62_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3376 U$$4335/A1 U$$3292/X _593_/Q U$$3293/X VGND VGND VPWR VPWR U$$3377/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2631 U$$28/A1 U$$2667/A2 U$$30/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2632/A sky130_fd_sc_hd__a22o_1
XU$$2642 U$$2642/A U$$2694/B VGND VGND VPWR VPWR U$$2642/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3387 U$$3387/A U$$3413/B VGND VGND VPWR VPWR U$$3387/X sky130_fd_sc_hd__xor2_1
XU$$2653 U$$50/A1 U$$2667/A2 U$$2790/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2654/A sky130_fd_sc_hd__a22o_1
XU$$3398 U$$4494/A1 U$$3292/X U$$4496/A1 U$$3293/X VGND VGND VPWR VPWR U$$3399/A sky130_fd_sc_hd__a22o_1
XFILLER_22_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2664 U$$2664/A U$$2710/B VGND VGND VPWR VPWR U$$2664/X sky130_fd_sc_hd__xor2_1
XU$$2675 _584_/Q U$$2607/X U$$4045/B1 U$$2608/X VGND VGND VPWR VPWR U$$2676/A sky130_fd_sc_hd__a22o_1
XU$$1930 U$$971/A1 U$$1922/X U$$12/B1 U$$1923/X VGND VGND VPWR VPWR U$$1931/A sky130_fd_sc_hd__a22o_1
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1941 U$$1941/A U$$1991/B VGND VGND VPWR VPWR U$$1941/X sky130_fd_sc_hd__xor2_1
XFILLER_34_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2686 U$$2686/A U$$2694/B VGND VGND VPWR VPWR U$$2686/X sky130_fd_sc_hd__xor2_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1952 U$$3457/B1 U$$2048/A2 U$$36/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1953/A sky130_fd_sc_hd__a22o_1
XU$$2697 U$$92/B1 U$$2729/A2 U$$96/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2698/A sky130_fd_sc_hd__a22o_1
XU$$1963 U$$1963/A U$$2023/B VGND VGND VPWR VPWR U$$1963/X sky130_fd_sc_hd__xor2_1
XU$$1974 U$$878/A1 U$$2036/A2 U$$880/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1975/A sky130_fd_sc_hd__a22o_1
XFILLER_15_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1985 U$$1985/A U$$1991/B VGND VGND VPWR VPWR U$$1985/X sky130_fd_sc_hd__xor2_1
XU$$1996 U$$78/A1 U$$2052/A2 U$$765/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$1997/A sky130_fd_sc_hd__a22o_1
XFILLER_193_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_98_0 dadda_fa_5_98_0/A dadda_fa_5_98_0/B dadda_fa_5_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/A dadda_fa_6_98_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_119_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$615 final_adder.U$$742/A final_adder.U$$742/B final_adder.U$$615/B1
+ VGND VGND VPWR VPWR final_adder.U$$743/B sky130_fd_sc_hd__a21o_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$626 final_adder.U$$626/A final_adder.U$$626/B VGND VGND VPWR VPWR
+ _172_/D sky130_fd_sc_hd__xor2_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$637 final_adder.U$$637/A final_adder.U$$637/B VGND VGND VPWR VPWR
+ _183_/D sky130_fd_sc_hd__xor2_1
XFILLER_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$648 final_adder.U$$648/A final_adder.U$$648/B VGND VGND VPWR VPWR
+ _194_/D sky130_fd_sc_hd__xor2_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$659 final_adder.U$$659/A final_adder.U$$659/B VGND VGND VPWR VPWR
+ _205_/D sky130_fd_sc_hd__xor2_1
XFILLER_99_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$509 U$$96/B1 U$$545/A2 U$$785/A1 U$$416/X VGND VGND VPWR VPWR U$$510/A sky130_fd_sc_hd__a22o_1
XU$$70 U$$70/A1 U$$4/X U$$70/B1 U$$5/X VGND VGND VPWR VPWR U$$71/A sky130_fd_sc_hd__a22o_1
XU$$81 U$$81/A U$$3/A VGND VGND VPWR VPWR U$$81/X sky130_fd_sc_hd__xor2_1
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$92 U$$92/A1 U$$4/X U$$92/B1 U$$5/X VGND VGND VPWR VPWR U$$93/A sky130_fd_sc_hd__a22o_1
XFILLER_72_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_107_1 U$$3812/X U$$3945/X U$$4078/X VGND VGND VPWR VPWR dadda_fa_4_108_0/CIN
+ dadda_fa_4_107_2/A sky130_fd_sc_hd__fa_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_48_3 dadda_fa_3_48_3/A dadda_fa_3_48_3/B dadda_fa_3_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/B dadda_fa_4_48_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1204 U$$928/B1 U$$1100/X _603_/Q U$$1101/X VGND VGND VPWR VPWR U$$1205/A sky130_fd_sc_hd__a22o_1
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1215 U$$1215/A U$$1232/A VGND VGND VPWR VPWR U$$1215/X sky130_fd_sc_hd__xor2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1226 U$$4514/A1 U$$1100/X _614_/Q U$$1101/X VGND VGND VPWR VPWR U$$1227/A sky130_fd_sc_hd__a22o_1
XFILLER_16_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1237 U$$1235/Y _634_/Q _633_/Q U$$1236/X U$$1233/Y VGND VGND VPWR VPWR U$$1237/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1248 U$$1248/A U$$1336/B VGND VGND VPWR VPWR U$$1248/X sky130_fd_sc_hd__xor2_1
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1259 _561_/Q U$$1341/A2 U$$987/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1260/A sky130_fd_sc_hd__a22o_1
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_50_3 dadda_fa_2_50_3/A dadda_fa_2_50_3/B dadda_fa_2_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/B dadda_fa_3_50_3/B sky130_fd_sc_hd__fa_2
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_43_2 U$$2753/X U$$2886/X input194/X VGND VGND VPWR VPWR dadda_fa_3_44_1/A
+ dadda_fa_3_43_3/A sky130_fd_sc_hd__fa_1
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3140 U$$4510/A1 U$$3146/A2 U$$950/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3141/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_20_1 dadda_fa_5_20_1/A dadda_fa_5_20_1/B dadda_fa_5_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/B dadda_fa_7_20_0/A sky130_fd_sc_hd__fa_1
XU$$3151 _661_/Q VGND VGND VPWR VPWR U$$3151/Y sky130_fd_sc_hd__inv_1
XU$$3162 U$$3162/A U$$3224/B VGND VGND VPWR VPWR U$$3162/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_1 U$$1143/X U$$1276/X U$$1409/X VGND VGND VPWR VPWR dadda_fa_3_37_0/CIN
+ dadda_fa_3_36_2/CIN sky130_fd_sc_hd__fa_1
XU$$3173 U$$979/B1 U$$3243/A2 U$$4271/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3174/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3184 U$$3184/A U$$3244/B VGND VGND VPWR VPWR U$$3184/X sky130_fd_sc_hd__xor2_1
XFILLER_35_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_13_0 dadda_fa_5_13_0/A dadda_fa_5_13_0/B dadda_fa_5_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/A dadda_fa_6_13_0/CIN sky130_fd_sc_hd__fa_1
XU$$2450 U$$2450/A U$$2464/B VGND VGND VPWR VPWR U$$2450/X sky130_fd_sc_hd__xor2_1
XU$$3195 U$$4291/A1 U$$3241/A2 U$$46/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3196/A sky130_fd_sc_hd__a22o_1
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_29_0 U$$65/X U$$198/X U$$331/X VGND VGND VPWR VPWR dadda_fa_3_30_1/B dadda_fa_3_29_3/A
+ sky130_fd_sc_hd__fa_2
XU$$2461 U$$4379/A1 U$$2463/A2 U$$956/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2462/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2472 U$$2472/A1 U$$2534/A2 U$$4255/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2473/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2483 U$$2483/A U$$2533/B VGND VGND VPWR VPWR U$$2483/X sky130_fd_sc_hd__xor2_1
XU$$2494 U$$28/A1 U$$2534/A2 U$$30/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2495/A sky130_fd_sc_hd__a22o_1
XFILLER_107_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1760 U$$938/A1 U$$1648/X U$$940/A1 U$$1649/X VGND VGND VPWR VPWR U$$1761/A sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1771 U$$1771/A _641_/Q VGND VGND VPWR VPWR U$$1771/X sky130_fd_sc_hd__xor2_1
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1782 _642_/Q VGND VGND VPWR VPWR U$$1784/B sky130_fd_sc_hd__inv_1
XU$$1793 U$$971/A1 U$$1867/A2 U$$12/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1794/A sky130_fd_sc_hd__a22o_1
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput70 b[14] VGND VGND VPWR VPWR _566_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput81 b[24] VGND VGND VPWR VPWR _576_/D sky130_fd_sc_hd__clkbuf_4
Xinput92 b[34] VGND VGND VPWR VPWR _586_/D sky130_fd_sc_hd__buf_2
XFILLER_190_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_58_2 dadda_fa_4_58_2/A dadda_fa_4_58_2/B dadda_fa_4_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/CIN dadda_fa_5_58_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$401 final_adder.U$$364/B final_adder.U$$718/B final_adder.U$$345/X
+ VGND VGND VPWR VPWR final_adder.U$$726/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$423 final_adder.U$$340/B final_adder.U$$702/B final_adder.U$$297/X
+ VGND VGND VPWR VPWR final_adder.U$$706/B sky130_fd_sc_hd__a21o_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$445 final_adder.U$$268/B final_adder.U$$646/B final_adder.U$$153/X
+ VGND VGND VPWR VPWR final_adder.U$$648/B sky130_fd_sc_hd__a21o_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_28_0 dadda_fa_7_28_0/A dadda_fa_7_28_0/B dadda_fa_7_28_0/CIN VGND VGND
+ VPWR VPWR _453_/D _324_/D sky130_fd_sc_hd__fa_2
Xrepeater660 _593_/Q VGND VGND VPWR VPWR U$$912/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$467 final_adder.U$$290/B final_adder.U$$690/B final_adder.U$$197/X
+ VGND VGND VPWR VPWR final_adder.U$$692/B sky130_fd_sc_hd__a21o_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater671 _589_/Q VGND VGND VPWR VPWR U$$630/A1 sky130_fd_sc_hd__buf_12
XU$$306 U$$32/A1 U$$278/X U$$34/A1 U$$279/X VGND VGND VPWR VPWR U$$307/A sky130_fd_sc_hd__a22o_1
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$317 U$$317/A U$$357/B VGND VGND VPWR VPWR U$$317/X sky130_fd_sc_hd__xor2_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater682 _585_/Q VGND VGND VPWR VPWR U$$4045/B1 sky130_fd_sc_hd__buf_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$489 final_adder.U$$312/B final_adder.U$$734/B final_adder.U$$241/X
+ VGND VGND VPWR VPWR final_adder.U$$736/B sky130_fd_sc_hd__a21o_1
XU$$328 U$$54/A1 U$$278/X U$$56/A1 U$$279/X VGND VGND VPWR VPWR U$$329/A sky130_fd_sc_hd__a22o_1
Xrepeater693 _581_/Q VGND VGND VPWR VPWR U$$3489/B1 sky130_fd_sc_hd__buf_12
XU$$339 U$$339/A U$$357/B VGND VGND VPWR VPWR U$$339/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_60_2 dadda_fa_3_60_2/A dadda_fa_3_60_2/B dadda_fa_3_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/A dadda_fa_4_60_2/B sky130_fd_sc_hd__fa_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_53_1 dadda_fa_3_53_1/A dadda_fa_3_53_1/B dadda_fa_3_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/CIN dadda_fa_4_53_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_69_1 U$$810/X U$$943/X U$$1076/X VGND VGND VPWR VPWR dadda_fa_1_70_6/B
+ dadda_fa_1_69_8/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_30_0 dadda_fa_6_30_0/A dadda_fa_6_30_0/B dadda_fa_6_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_31_0/B dadda_fa_7_30_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_46_0 dadda_fa_3_46_0/A dadda_fa_3_46_0/B dadda_fa_3_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/B dadda_fa_4_46_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$840 U$$18/A1 U$$928/A2 U$$842/A1 U$$928/B2 VGND VGND VPWR VPWR U$$841/A sky130_fd_sc_hd__a22o_1
X_677_ _677_/CLK _677_/D VGND VGND VPWR VPWR _677_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$851 U$$851/A U$$923/B VGND VGND VPWR VPWR U$$851/X sky130_fd_sc_hd__xor2_1
XU$$862 U$$40/A1 U$$928/A2 _569_/Q U$$928/B2 VGND VGND VPWR VPWR U$$863/A sky130_fd_sc_hd__a22o_1
XU$$1001 U$$3876/B1 U$$999/A2 U$$4291/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1002/A sky130_fd_sc_hd__a22o_1
XU$$1012 U$$1012/A U$$980/B VGND VGND VPWR VPWR U$$1012/X sky130_fd_sc_hd__xor2_1
XU$$873 U$$873/A U$$903/B VGND VGND VPWR VPWR U$$873/X sky130_fd_sc_hd__xor2_1
XU$$884 U$$62/A1 U$$910/A2 U$$64/A1 U$$910/B2 VGND VGND VPWR VPWR U$$885/A sky130_fd_sc_hd__a22o_1
XU$$1023 U$$64/A1 U$$999/A2 U$$66/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1024/A sky130_fd_sc_hd__a22o_1
XU$$1034 U$$1034/A U$$980/B VGND VGND VPWR VPWR U$$1034/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$895 U$$895/A U$$903/B VGND VGND VPWR VPWR U$$895/X sky130_fd_sc_hd__xor2_1
XU$$1045 U$$908/A1 U$$1093/A2 U$$88/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1046/A sky130_fd_sc_hd__a22o_1
XU$$1056 U$$1056/A U$$998/B VGND VGND VPWR VPWR U$$1056/X sky130_fd_sc_hd__xor2_1
XFILLER_188_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1067 U$$930/A1 U$$963/X U$$932/A1 U$$964/X VGND VGND VPWR VPWR U$$1068/A sky130_fd_sc_hd__a22o_1
XU$$1078 U$$1078/A U$$998/B VGND VGND VPWR VPWR U$$1078/X sky130_fd_sc_hd__xor2_1
XU$$1089 U$$952/A1 U$$963/X U$$952/B1 U$$964/X VGND VGND VPWR VPWR U$$1090/A sky130_fd_sc_hd__a22o_1
XFILLER_176_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_103_0 dadda_fa_7_103_0/A dadda_fa_7_103_0/B dadda_fa_7_103_0/CIN VGND
+ VGND VPWR VPWR _528_/D _399_/D sky130_fd_sc_hd__fa_2
XFILLER_129_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_98_3 U$$3528/X U$$3661/X U$$3794/X VGND VGND VPWR VPWR dadda_fa_3_99_1/CIN
+ dadda_fa_3_98_3/B sky130_fd_sc_hd__fa_1
XFILLER_176_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_688__908 VGND VGND VPWR VPWR _688__908/HI _688__908/LO sky130_fd_sc_hd__conb_1
XFILLER_171_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_68_1 dadda_fa_5_68_1/A dadda_fa_5_68_1/B dadda_fa_5_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/B dadda_fa_7_68_0/A sky130_fd_sc_hd__fa_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_107_0 U$$3013/Y U$$3147/X U$$3280/X VGND VGND VPWR VPWR dadda_fa_3_108_3/CIN
+ dadda_fa_4_107_0/A sky130_fd_sc_hd__fa_1
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2280 U$$4335/A1 U$$2326/A2 _593_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2281/A sky130_fd_sc_hd__a22o_1
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2291 U$$2291/A U$$2327/B VGND VGND VPWR VPWR U$$2291/X sky130_fd_sc_hd__xor2_1
XFILLER_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1590 U$$1590/A U$$1614/B VGND VGND VPWR VPWR U$$1590/X sky130_fd_sc_hd__xor2_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_70_1 dadda_fa_4_70_1/A dadda_fa_4_70_1/B dadda_fa_4_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/B dadda_fa_5_70_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_1 U$$1908/X U$$2041/X U$$2174/X VGND VGND VPWR VPWR dadda_fa_2_87_3/A
+ dadda_fa_2_86_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_63_0 dadda_fa_4_63_0/A dadda_fa_4_63_0/B dadda_fa_4_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/A dadda_fa_5_63_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_0 U$$1095/Y U$$1229/X U$$1362/X VGND VGND VPWR VPWR dadda_fa_2_80_0/B
+ dadda_fa_2_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$220 final_adder.U$$715/A final_adder.U$$714/A VGND VGND VPWR VPWR
+ final_adder.U$$302/B sky130_fd_sc_hd__and2_1
XFILLER_131_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$231 final_adder.U$$725/A final_adder.U$$597/B1 final_adder.U$$231/B1
+ VGND VGND VPWR VPWR final_adder.U$$231/X sky130_fd_sc_hd__a21o_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$242 final_adder.U$$737/A final_adder.U$$736/A VGND VGND VPWR VPWR
+ final_adder.U$$312/A sky130_fd_sc_hd__and2_1
X_600_ _601_/CLK _600_/D VGND VGND VPWR VPWR _600_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3909 U$$3909/A U$$3929/B VGND VGND VPWR VPWR U$$3909/X sky130_fd_sc_hd__xor2_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$253 final_adder.U$$747/A final_adder.U$$619/B1 final_adder.U$$253/B1
+ VGND VGND VPWR VPWR final_adder.U$$253/X sky130_fd_sc_hd__a21o_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$264 final_adder.U$$264/A final_adder.U$$264/B VGND VGND VPWR VPWR
+ final_adder.U$$324/B sky130_fd_sc_hd__and2_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$103 U$$103/A U$$3/A VGND VGND VPWR VPWR U$$103/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$275 final_adder.U$$274/A final_adder.U$$165/X final_adder.U$$167/X
+ VGND VGND VPWR VPWR final_adder.U$$275/X sky130_fd_sc_hd__a21o_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$114 U$$799/A1 U$$4/X U$$938/A1 U$$5/X VGND VGND VPWR VPWR U$$115/A sky130_fd_sc_hd__a22o_1
XFILLER_73_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$286 final_adder.U$$286/A final_adder.U$$286/B VGND VGND VPWR VPWR
+ final_adder.U$$334/A sky130_fd_sc_hd__and2_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$125 U$$125/A U$$3/A VGND VGND VPWR VPWR U$$125/X sky130_fd_sc_hd__xor2_1
Xrepeater490 U$$2334/X VGND VGND VPWR VPWR U$$2463/B2 sky130_fd_sc_hd__buf_12
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_531_ _531_/CLK _531_/D VGND VGND VPWR VPWR _531_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$297 final_adder.U$$296/A final_adder.U$$209/X final_adder.U$$211/X
+ VGND VGND VPWR VPWR final_adder.U$$297/X sky130_fd_sc_hd__a21o_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$136 U$$89/B VGND VGND VPWR VPWR U$$136/Y sky130_fd_sc_hd__inv_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$147 U$$8/B1 U$$141/X U$$12/A1 U$$142/X VGND VGND VPWR VPWR U$$148/A sky130_fd_sc_hd__a22o_1
XFILLER_26_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$158 U$$158/A U$$274/A VGND VGND VPWR VPWR U$$158/X sky130_fd_sc_hd__xor2_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$169 U$$32/A1 U$$141/X U$$34/A1 U$$142/X VGND VGND VPWR VPWR U$$170/A sky130_fd_sc_hd__a22o_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ _462_/CLK _462_/D VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_393_ _595_/CLK _393_/D VGND VGND VPWR VPWR _393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_78_0 dadda_fa_6_78_0/A dadda_fa_6_78_0/B dadda_fa_6_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_79_0/B dadda_fa_7_78_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$670 U$$944/A1 U$$552/X U$$946/A1 U$$553/X VGND VGND VPWR VPWR U$$671/A sky130_fd_sc_hd__a22o_1
XU$$681 U$$681/A _625_/Q VGND VGND VPWR VPWR U$$681/X sky130_fd_sc_hd__xor2_1
XFILLER_32_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$692 U$$692/A U$$784/B VGND VGND VPWR VPWR U$$692/X sky130_fd_sc_hd__xor2_1
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_770__822 VGND VGND VPWR VPWR _770__822/HI U$$4388/A2 sky130_fd_sc_hd__conb_1
XFILLER_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_80_0 dadda_fa_5_80_0/A dadda_fa_5_80_0/B dadda_fa_5_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/A dadda_fa_6_80_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_96_0 U$$2460/X U$$2593/X U$$2726/X VGND VGND VPWR VPWR dadda_fa_3_97_0/B
+ dadda_fa_3_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_811__863 VGND VGND VPWR VPWR _811__863/HI U$$4467/B sky130_fd_sc_hd__conb_1
XFILLER_87_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_72_7 dadda_fa_1_72_7/A dadda_fa_1_72_7/B dadda_fa_1_72_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_2/CIN dadda_fa_2_72_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_65_6 dadda_fa_1_65_6/A dadda_fa_1_65_6/B dadda_fa_1_65_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/B dadda_fa_2_65_5/B sky130_fd_sc_hd__fa_1
XFILLER_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_58_5 U$$3581/X U$$3714/X U$$3847/X VGND VGND VPWR VPWR dadda_fa_2_59_2/A
+ dadda_fa_2_58_5/A sky130_fd_sc_hd__fa_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_95_0 dadda_fa_7_95_0/A dadda_fa_7_95_0/B dadda_fa_7_95_0/CIN VGND VGND
+ VPWR VPWR _520_/D _391_/D sky130_fd_sc_hd__fa_2
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4407 U$$4407/A U$$4407/B VGND VGND VPWR VPWR U$$4407/X sky130_fd_sc_hd__xor2_2
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4418 _565_/Q U$$4388/X _566_/Q U$$4389/X VGND VGND VPWR VPWR U$$4419/A sky130_fd_sc_hd__a22o_1
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4429 U$$4429/A U$$4429/B VGND VGND VPWR VPWR U$$4429/X sky130_fd_sc_hd__xor2_2
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_110_0 dadda_fa_6_110_0/A dadda_fa_6_110_0/B dadda_fa_6_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_111_0/B dadda_fa_7_110_0/CIN sky130_fd_sc_hd__fa_2
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3706 U$$3706/A U$$3756/B VGND VGND VPWR VPWR U$$3706/X sky130_fd_sc_hd__xor2_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3717 U$$975/B1 U$$3795/A2 U$$979/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3718/A sky130_fd_sc_hd__a22o_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3728 U$$3728/A U$$3784/B VGND VGND VPWR VPWR U$$3728/X sky130_fd_sc_hd__xor2_1
XU$$3739 U$$4424/A1 U$$3795/A2 U$$4289/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3740/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_3 dadda_fa_3_30_3/A dadda_fa_3_30_3/B dadda_fa_3_30_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/B dadda_fa_4_30_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_514_ _518_/CLK _514_/D VGND VGND VPWR VPWR _514_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_3_23_2 U$$1117/X U$$1250/X U$$1383/X VGND VGND VPWR VPWR dadda_fa_4_24_1/A
+ dadda_fa_4_23_2/B sky130_fd_sc_hd__fa_1
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_445_ _461_/CLK _445_/D VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _509_/CLK _376_/D VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_754__806 VGND VGND VPWR VPWR _754__806/HI U$$3705/A1 sky130_fd_sc_hd__conb_1
XFILLER_174_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_75_5 dadda_fa_2_75_5/A dadda_fa_2_75_5/B dadda_fa_2_75_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_2/A dadda_fa_4_75_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_4 dadda_fa_2_68_4/A dadda_fa_2_68_4/B dadda_fa_2_68_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/CIN dadda_fa_3_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_105_1 dadda_fa_5_105_1/A dadda_fa_5_105_1/B dadda_fa_5_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/B dadda_fa_7_105_0/A sky130_fd_sc_hd__fa_2
XFILLER_173_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_70_4 U$$3871/X U$$4004/X U$$4137/X VGND VGND VPWR VPWR dadda_fa_2_71_1/CIN
+ dadda_fa_2_70_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_63_3 U$$3591/X U$$3724/X U$$3857/X VGND VGND VPWR VPWR dadda_fa_2_64_1/B
+ dadda_fa_2_63_4/B sky130_fd_sc_hd__fa_2
XFILLER_75_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_40_2 dadda_fa_4_40_2/A dadda_fa_4_40_2/B dadda_fa_4_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/CIN dadda_fa_5_40_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_189_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_56_2 U$$1981/X U$$2114/X U$$2247/X VGND VGND VPWR VPWR dadda_fa_2_57_1/A
+ dadda_fa_2_56_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_33_1 dadda_fa_4_33_1/A dadda_fa_4_33_1/B dadda_fa_4_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/B dadda_fa_5_33_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_1 U$$504/X U$$637/X U$$770/X VGND VGND VPWR VPWR dadda_fa_2_50_1/A
+ dadda_fa_2_49_4/A sky130_fd_sc_hd__fa_2
XFILLER_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_10_0 dadda_fa_7_10_0/A dadda_fa_7_10_0/B dadda_fa_7_10_0/CIN VGND VGND
+ VPWR VPWR _435_/D _306_/D sky130_fd_sc_hd__fa_2
XFILLER_43_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_26_0 dadda_fa_4_26_0/A dadda_fa_4_26_0/B dadda_fa_4_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/A dadda_fa_5_26_1/A sky130_fd_sc_hd__fa_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_230_ _499_/CLK _230_/D VGND VGND VPWR VPWR _230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_78_3 dadda_fa_3_78_3/A dadda_fa_3_78_3/B dadda_fa_3_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/B dadda_fa_4_78_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4204 U$$94/A1 U$$4244/A2 U$$94/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4205/A sky130_fd_sc_hd__a22o_1
XFILLER_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4215 U$$4215/A U$$4246/A VGND VGND VPWR VPWR U$$4215/X sky130_fd_sc_hd__xor2_1
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4226 U$$4500/A1 U$$4244/A2 U$$4502/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4227/A
+ sky130_fd_sc_hd__a22o_1
XU$$4237 U$$4237/A U$$4246/A VGND VGND VPWR VPWR U$$4237/X sky130_fd_sc_hd__xor2_1
XFILLER_120_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_3_15_0 U$$37/X U$$170/X VGND VGND VPWR VPWR dadda_fa_4_16_2/A dadda_ha_3_15_0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3503 U$$78/A1 U$$3545/A2 U$$765/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3504/A sky130_fd_sc_hd__a22o_1
XU$$4248 _678_/Q VGND VGND VPWR VPWR U$$4250/B sky130_fd_sc_hd__inv_1
XU$$3514 U$$3514/A U$$3536/B VGND VGND VPWR VPWR U$$3514/X sky130_fd_sc_hd__xor2_1
XU$$4259 _554_/Q U$$4381/A2 _555_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4260/A sky130_fd_sc_hd__a22o_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3525 U$$4484/A1 U$$3525/A2 _599_/Q U$$3525/B2 VGND VGND VPWR VPWR U$$3526/A sky130_fd_sc_hd__a22o_1
XU$$3536 U$$3536/A U$$3536/B VGND VGND VPWR VPWR U$$3536/X sky130_fd_sc_hd__xor2_1
XFILLER_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2802 U$$3624/A1 U$$2868/A2 U$$3900/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2803/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3547 U$$4506/A1 U$$3429/X U$$4508/A1 U$$3430/X VGND VGND VPWR VPWR U$$3548/A sky130_fd_sc_hd__a22o_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2813 U$$2813/A U$$2871/B VGND VGND VPWR VPWR U$$2813/X sky130_fd_sc_hd__xor2_1
XU$$3558 U$$3558/A U$$3561/A VGND VGND VPWR VPWR U$$3558/X sky130_fd_sc_hd__xor2_1
XFILLER_18_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3569 U$$3569/A U$$3698/A VGND VGND VPWR VPWR U$$3569/X sky130_fd_sc_hd__xor2_1
XFILLER_46_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2824 U$$632/A1 U$$2868/A2 U$$771/A1 U$$2745/X VGND VGND VPWR VPWR U$$2825/A sky130_fd_sc_hd__a22o_1
XU$$2835 U$$2835/A U$$2871/B VGND VGND VPWR VPWR U$$2835/X sky130_fd_sc_hd__xor2_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2846 _601_/Q U$$2868/A2 U$$928/B1 U$$2870/B2 VGND VGND VPWR VPWR U$$2847/A sky130_fd_sc_hd__a22o_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2857 U$$2857/A U$$2871/B VGND VGND VPWR VPWR U$$2857/X sky130_fd_sc_hd__xor2_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2868 U$$950/A1 U$$2868/A2 U$$4514/A1 U$$2870/B2 VGND VGND VPWR VPWR U$$2869/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2879 _659_/Q VGND VGND VPWR VPWR U$$2879/Y sky130_fd_sc_hd__inv_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _432_/CLK _428_/D VGND VGND VPWR VPWR _428_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_359_ _488_/CLK _359_/D VGND VGND VPWR VPWR _359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_80_3 dadda_fa_2_80_3/A dadda_fa_2_80_3/B dadda_fa_2_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/B dadda_fa_3_80_3/B sky130_fd_sc_hd__fa_2
XFILLER_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_73_2 dadda_fa_2_73_2/A dadda_fa_2_73_2/B dadda_fa_2_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/A dadda_fa_3_73_3/A sky130_fd_sc_hd__fa_2
Xdadda_fa_5_50_1 dadda_fa_5_50_1/A dadda_fa_5_50_1/B dadda_fa_5_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/B dadda_fa_7_50_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_66_1 dadda_fa_2_66_1/A dadda_fa_2_66_1/B dadda_fa_2_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/CIN dadda_fa_3_66_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_43_0 dadda_fa_5_43_0/A dadda_fa_5_43_0/B dadda_fa_5_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/A dadda_fa_6_43_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_59_0 dadda_fa_2_59_0/A dadda_fa_2_59_0/B dadda_fa_2_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/B dadda_fa_3_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput2 a[10] VGND VGND VPWR VPWR _626_/D sky130_fd_sc_hd__buf_2
XFILLER_7_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$0 _424_/Q _296_/Q VGND VGND VPWR VPWR final_adder.U$$623/B final_adder.U$$622/A
+ sky130_fd_sc_hd__ha_1
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_88_2 dadda_fa_4_88_2/A dadda_fa_4_88_2/B dadda_fa_4_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/CIN dadda_fa_5_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput350 _237_/Q VGND VGND VPWR VPWR o[69] sky130_fd_sc_hd__buf_2
XFILLER_156_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput361 _247_/Q VGND VGND VPWR VPWR o[79] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_58_0 dadda_fa_7_58_0/A dadda_fa_7_58_0/B dadda_fa_7_58_0/CIN VGND VGND
+ VPWR VPWR _483_/D _354_/D sky130_fd_sc_hd__fa_1
Xoutput372 _257_/Q VGND VGND VPWR VPWR o[89] sky130_fd_sc_hd__buf_2
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput383 _267_/Q VGND VGND VPWR VPWR o[99] sky130_fd_sc_hd__buf_2
XFILLER_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_61_0 U$$1991/X U$$2124/X U$$2257/X VGND VGND VPWR VPWR dadda_fa_2_62_0/B
+ dadda_fa_2_61_3/B sky130_fd_sc_hd__fa_2
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2109 U$$4438/A1 U$$2117/A2 U$$878/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2110/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1408 U$$38/A1 U$$1474/A2 U$$3191/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1409/A sky130_fd_sc_hd__a22o_1
XU$$1419 U$$1419/A U$$1461/B VGND VGND VPWR VPWR U$$1419/X sky130_fd_sc_hd__xor2_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ _480_/CLK _213_/D VGND VGND VPWR VPWR _213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_90_2 dadda_fa_3_90_2/A dadda_fa_3_90_2/B dadda_fa_3_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/A dadda_fa_4_90_2/B sky130_fd_sc_hd__fa_1
XFILLER_125_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_83_1 dadda_fa_3_83_1/A dadda_fa_3_83_1/B dadda_fa_3_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/CIN dadda_fa_4_83_2/A sky130_fd_sc_hd__fa_2
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_60_0 dadda_fa_6_60_0/A dadda_fa_6_60_0/B dadda_fa_6_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_61_0/B dadda_fa_7_60_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_76_0 dadda_fa_3_76_0/A dadda_fa_3_76_0/B dadda_fa_3_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/B dadda_fa_4_76_1/CIN sky130_fd_sc_hd__fa_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4001 _562_/Q U$$3977/X _563_/Q U$$3978/X VGND VGND VPWR VPWR U$$4002/A sky130_fd_sc_hd__a22o_1
XU$$4012 U$$4012/A U$$4109/A VGND VGND VPWR VPWR U$$4012/X sky130_fd_sc_hd__xor2_1
XFILLER_93_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4023 _573_/Q U$$3977/X U$$50/B1 U$$3978/X VGND VGND VPWR VPWR U$$4024/A sky130_fd_sc_hd__a22o_1
XFILLER_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4034 U$$4034/A U$$4044/B VGND VGND VPWR VPWR U$$4034/X sky130_fd_sc_hd__xor2_1
XU$$4045 _584_/Q U$$4045/A2 U$$4045/B1 U$$3978/X VGND VGND VPWR VPWR U$$4046/A sky130_fd_sc_hd__a22o_1
XU$$3300 U$$4122/A1 U$$3396/A2 U$$14/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3301/A sky130_fd_sc_hd__a22o_1
XU$$3311 U$$3311/A U$$3413/B VGND VGND VPWR VPWR U$$3311/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_1 dadda_fa_4_112_1/A dadda_fa_4_112_1/B dadda_fa_4_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/B dadda_fa_5_112_1/B sky130_fd_sc_hd__fa_1
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4056 U$$4056/A U$$4058/B VGND VGND VPWR VPWR U$$4056/X sky130_fd_sc_hd__xor2_1
XU$$4067 U$$94/A1 U$$4107/A2 _596_/Q U$$4107/B2 VGND VGND VPWR VPWR U$$4068/A sky130_fd_sc_hd__a22o_1
XU$$3322 U$$3457/B1 U$$3396/A2 U$$4283/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3323/A
+ sky130_fd_sc_hd__a22o_1
XU$$4078 U$$4078/A _675_/Q VGND VGND VPWR VPWR U$$4078/X sky130_fd_sc_hd__xor2_1
XU$$3333 U$$3333/A U$$3413/B VGND VGND VPWR VPWR U$$3333/X sky130_fd_sc_hd__xor2_1
XU$$3344 U$$4303/A1 U$$3292/X _577_/Q U$$3293/X VGND VGND VPWR VPWR U$$3345/A sky130_fd_sc_hd__a22o_1
XU$$4089 U$$4500/A1 U$$4107/A2 U$$4502/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4090/A
+ sky130_fd_sc_hd__a22o_1
XU$$3355 U$$3355/A U$$3403/B VGND VGND VPWR VPWR U$$3355/X sky130_fd_sc_hd__xor2_1
XFILLER_47_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2610 U$$2610/A U$$2710/B VGND VGND VPWR VPWR U$$2610/X sky130_fd_sc_hd__xor2_1
XU$$2621 U$$4265/A1 U$$2667/A2 U$$979/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2622/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_105_0 dadda_fa_4_105_0/A dadda_fa_4_105_0/B dadda_fa_4_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/A dadda_fa_5_105_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_38_5 dadda_fa_2_38_5/A dadda_fa_2_38_5/B dadda_fa_2_38_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_39_2/A dadda_fa_4_38_0/A sky130_fd_sc_hd__fa_2
XU$$3366 _587_/Q U$$3292/X _588_/Q U$$3293/X VGND VGND VPWR VPWR U$$3367/A sky130_fd_sc_hd__a22o_1
XU$$3377 U$$3377/A U$$3403/B VGND VGND VPWR VPWR U$$3377/X sky130_fd_sc_hd__xor2_1
XU$$2632 U$$2632/A U$$2694/B VGND VGND VPWR VPWR U$$2632/X sky130_fd_sc_hd__xor2_1
XU$$2643 U$$3191/A1 U$$2667/A2 U$$4289/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2644/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3388 U$$4484/A1 U$$3292/X _599_/Q U$$3293/X VGND VGND VPWR VPWR U$$3389/A sky130_fd_sc_hd__a22o_1
XU$$3399 U$$3399/A U$$3403/B VGND VGND VPWR VPWR U$$3399/X sky130_fd_sc_hd__xor2_1
XU$$2654 U$$2654/A U$$2694/B VGND VGND VPWR VPWR U$$2654/X sky130_fd_sc_hd__xor2_1
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1920 U$$2055/A VGND VGND VPWR VPWR U$$1920/Y sky130_fd_sc_hd__inv_1
XFILLER_55_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2665 U$$4446/A1 U$$2729/A2 U$$64/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2666/A sky130_fd_sc_hd__a22o_1
XU$$2676 U$$2676/A U$$2698/B VGND VGND VPWR VPWR U$$2676/X sky130_fd_sc_hd__xor2_1
XU$$1931 U$$1931/A U$$2021/B VGND VGND VPWR VPWR U$$1931/X sky130_fd_sc_hd__xor2_1
XU$$1942 U$$983/A1 U$$1922/X U$$26/A1 U$$1923/X VGND VGND VPWR VPWR U$$1943/A sky130_fd_sc_hd__a22o_1
XFILLER_61_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2687 _590_/Q U$$2607/X _591_/Q U$$2608/X VGND VGND VPWR VPWR U$$2688/A sky130_fd_sc_hd__a22o_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2698 U$$2698/A U$$2698/B VGND VGND VPWR VPWR U$$2698/X sky130_fd_sc_hd__xor2_1
XU$$1953 U$$1953/A U$$1991/B VGND VGND VPWR VPWR U$$1953/X sky130_fd_sc_hd__xor2_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1964 U$$868/A1 U$$1922/X U$$48/A1 U$$1923/X VGND VGND VPWR VPWR U$$1965/A sky130_fd_sc_hd__a22o_1
XU$$1975 U$$1975/A U$$1991/B VGND VGND VPWR VPWR U$$1975/X sky130_fd_sc_hd__xor2_1
XU$$1986 U$$3217/B1 U$$2036/A2 U$$892/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1987/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1997 U$$1997/A U$$2021/B VGND VGND VPWR VPWR U$$1997/X sky130_fd_sc_hd__xor2_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_98_1 dadda_fa_5_98_1/A dadda_fa_5_98_1/B dadda_fa_5_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/B dadda_fa_7_98_0/A sky130_fd_sc_hd__fa_2
XFILLER_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$605 final_adder.U$$732/A final_adder.U$$732/B final_adder.U$$605/B1
+ VGND VGND VPWR VPWR final_adder.U$$733/B sky130_fd_sc_hd__a21o_1
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$627 final_adder.U$$627/A final_adder.U$$627/B VGND VGND VPWR VPWR
+ _173_/D sky130_fd_sc_hd__xor2_2
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$638 final_adder.U$$638/A final_adder.U$$638/B VGND VGND VPWR VPWR
+ _184_/D sky130_fd_sc_hd__xor2_1
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$649 final_adder.U$$649/A final_adder.U$$649/B VGND VGND VPWR VPWR
+ _195_/D sky130_fd_sc_hd__xor2_2
XFILLER_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$60 U$$60/A1 U$$4/X U$$62/A1 U$$5/X VGND VGND VPWR VPWR U$$61/A sky130_fd_sc_hd__a22o_1
XU$$71 U$$71/A U$$89/B VGND VGND VPWR VPWR U$$71/X sky130_fd_sc_hd__xor2_1
XFILLER_65_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$82 U$$82/A1 U$$4/X U$$84/A1 U$$5/X VGND VGND VPWR VPWR U$$83/A sky130_fd_sc_hd__a22o_1
XU$$93 U$$93/A U$$3/A VGND VGND VPWR VPWR U$$93/X sky130_fd_sc_hd__xor2_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_93_0 dadda_fa_4_93_0/A dadda_fa_4_93_0/B dadda_fa_4_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/A dadda_fa_5_93_1/A sky130_fd_sc_hd__fa_1
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_2 U$$4211/X U$$4344/X U$$4477/X VGND VGND VPWR VPWR dadda_fa_4_108_1/A
+ dadda_fa_4_107_2/B sky130_fd_sc_hd__fa_2
XFILLER_134_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1205 U$$1205/A U$$1232/A VGND VGND VPWR VPWR U$$1205/X sky130_fd_sc_hd__xor2_1
XU$$1216 U$$4504/A1 U$$1100/X U$$944/A1 U$$1101/X VGND VGND VPWR VPWR U$$1217/A sky130_fd_sc_hd__a22o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1227 U$$1227/A U$$1232/A VGND VGND VPWR VPWR U$$1227/X sky130_fd_sc_hd__xor2_1
XU$$1238 U$$1236/B _633_/Q _634_/Q U$$1233/Y VGND VGND VPWR VPWR U$$1238/X sky130_fd_sc_hd__a22o_4
XU$$1249 U$$14/B1 U$$1237/X U$$18/A1 U$$1238/X VGND VGND VPWR VPWR U$$1250/A sky130_fd_sc_hd__a22o_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_50_4 dadda_fa_2_50_4/A dadda_fa_2_50_4/B dadda_fa_2_50_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/CIN dadda_fa_3_50_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_43_3 dadda_fa_2_43_3/A dadda_fa_2_43_3/B dadda_fa_2_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/B dadda_fa_3_43_3/B sky130_fd_sc_hd__fa_1
XFILLER_94_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3130 _606_/Q U$$3018/X _607_/Q U$$3019/X VGND VGND VPWR VPWR U$$3131/A sky130_fd_sc_hd__a22o_1
XFILLER_47_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3141 U$$3141/A _661_/Q VGND VGND VPWR VPWR U$$3141/X sky130_fd_sc_hd__xor2_1
XU$$3152 _662_/Q VGND VGND VPWR VPWR U$$3154/B sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_2 U$$1542/X U$$1675/X U$$1808/X VGND VGND VPWR VPWR dadda_fa_3_37_1/A
+ dadda_fa_3_36_3/A sky130_fd_sc_hd__fa_2
XU$$3163 U$$12/A1 U$$3241/A2 _555_/Q U$$3253/B2 VGND VGND VPWR VPWR U$$3164/A sky130_fd_sc_hd__a22o_1
XU$$3174 U$$3174/A U$$3244/B VGND VGND VPWR VPWR U$$3174/X sky130_fd_sc_hd__xor2_2
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2440 U$$2440/A U$$2464/B VGND VGND VPWR VPWR U$$2440/X sky130_fd_sc_hd__xor2_1
XU$$3185 U$$3457/B1 U$$3241/A2 U$$4283/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3186/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_13_1 dadda_fa_5_13_1/A dadda_fa_5_13_1/B dadda_ha_4_13_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/B dadda_fa_7_13_0/A sky130_fd_sc_hd__fa_2
XFILLER_185_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_29_1 U$$464/X U$$597/X U$$730/X VGND VGND VPWR VPWR dadda_fa_3_30_1/CIN
+ dadda_fa_3_29_3/B sky130_fd_sc_hd__fa_1
XU$$3196 U$$3196/A U$$3224/B VGND VGND VPWR VPWR U$$3196/X sky130_fd_sc_hd__xor2_1
XU$$2451 _609_/Q U$$2463/A2 _610_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2452/A sky130_fd_sc_hd__a22o_1
XU$$2462 U$$2462/A U$$2464/B VGND VGND VPWR VPWR U$$2462/X sky130_fd_sc_hd__xor2_1
XU$$2473 U$$2473/A U$$2533/B VGND VGND VPWR VPWR U$$2473/X sky130_fd_sc_hd__xor2_2
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2484 U$$4265/A1 U$$2534/A2 U$$979/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2485/A
+ sky130_fd_sc_hd__a22o_1
XU$$1750 U$$928/A1 U$$1770/A2 _602_/Q U$$1770/B2 VGND VGND VPWR VPWR U$$1751/A sky130_fd_sc_hd__a22o_1
XU$$2495 U$$2495/A U$$2585/B VGND VGND VPWR VPWR U$$2495/X sky130_fd_sc_hd__xor2_1
XU$$1761 U$$1761/A U$$1781/A VGND VGND VPWR VPWR U$$1761/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1772 U$$950/A1 U$$1648/X U$$4514/A1 U$$1649/X VGND VGND VPWR VPWR U$$1773/A sky130_fd_sc_hd__a22o_1
XU$$1783 U$$1918/A VGND VGND VPWR VPWR U$$1783/Y sky130_fd_sc_hd__inv_1
XU$$1794 U$$1794/A U$$1918/A VGND VGND VPWR VPWR U$$1794/X sky130_fd_sc_hd__xor2_1
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput60 a[63] VGND VGND VPWR VPWR _679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput71 b[15] VGND VGND VPWR VPWR _567_/D sky130_fd_sc_hd__clkbuf_4
Xinput82 b[25] VGND VGND VPWR VPWR _577_/D sky130_fd_sc_hd__clkbuf_4
Xinput93 b[35] VGND VGND VPWR VPWR _587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$413 final_adder.U$$330/B final_adder.U$$662/B final_adder.U$$277/X
+ VGND VGND VPWR VPWR final_adder.U$$666/B sky130_fd_sc_hd__a21o_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$435 final_adder.U$$258/B final_adder.U$$626/B final_adder.U$$133/X
+ VGND VGND VPWR VPWR final_adder.U$$628/B sky130_fd_sc_hd__a21o_1
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater650 _597_/Q VGND VGND VPWR VPWR U$$98/A1 sky130_fd_sc_hd__buf_12
XFILLER_96_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$457 final_adder.U$$280/B final_adder.U$$670/B final_adder.U$$177/X
+ VGND VGND VPWR VPWR final_adder.U$$672/B sky130_fd_sc_hd__a21o_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater661 U$$771/B1 VGND VGND VPWR VPWR U$$88/A1 sky130_fd_sc_hd__buf_12
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$307 U$$307/A U$$357/B VGND VGND VPWR VPWR U$$307/X sky130_fd_sc_hd__xor2_1
Xrepeater672 _588_/Q VGND VGND VPWR VPWR U$$902/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$479 final_adder.U$$302/B final_adder.U$$714/B final_adder.U$$221/X
+ VGND VGND VPWR VPWR final_adder.U$$716/B sky130_fd_sc_hd__a21o_1
XU$$318 _570_/Q U$$278/X U$$46/A1 U$$279/X VGND VGND VPWR VPWR U$$319/A sky130_fd_sc_hd__a22o_1
Xrepeater683 U$$72/A1 VGND VGND VPWR VPWR U$$70/B1 sky130_fd_sc_hd__buf_12
XU$$329 U$$329/A U$$391/B VGND VGND VPWR VPWR U$$329/X sky130_fd_sc_hd__xor2_1
Xrepeater694 _580_/Q VGND VGND VPWR VPWR U$$64/A1 sky130_fd_sc_hd__buf_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_112_0 _699__919/HI U$$3423/X U$$3556/X VGND VGND VPWR VPWR dadda_fa_4_113_1/B
+ dadda_fa_4_112_2/A sky130_fd_sc_hd__fa_1
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_60_3 dadda_fa_3_60_3/A dadda_fa_3_60_3/B dadda_fa_3_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/B dadda_fa_4_60_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_53_2 dadda_fa_3_53_2/A dadda_fa_3_53_2/B dadda_fa_3_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/A dadda_fa_4_53_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_69_2 U$$1209/X U$$1342/X U$$1475/X VGND VGND VPWR VPWR dadda_fa_1_70_6/CIN
+ dadda_fa_1_69_8/B sky130_fd_sc_hd__fa_1
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_46_1 dadda_fa_3_46_1/A dadda_fa_3_46_1/B dadda_fa_3_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/CIN dadda_fa_4_46_2/A sky130_fd_sc_hd__fa_1
XFILLER_17_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_23_0 dadda_fa_6_23_0/A dadda_fa_6_23_0/B dadda_fa_6_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_24_0/B dadda_fa_7_23_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_17_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_39_0 dadda_fa_3_39_0/A dadda_fa_3_39_0/B dadda_fa_3_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/B dadda_fa_4_39_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_21_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$830 U$$8/A1 U$$928/A2 U$$8/B1 U$$928/B2 VGND VGND VPWR VPWR U$$831/A sky130_fd_sc_hd__a22o_1
X_676_ _678_/CLK _676_/D VGND VGND VPWR VPWR _676_/Q sky130_fd_sc_hd__dfxtp_1
XU$$841 U$$841/A U$$923/B VGND VGND VPWR VPWR U$$841/X sky130_fd_sc_hd__xor2_1
XU$$852 U$$28/B1 U$$910/A2 U$$32/A1 U$$910/B2 VGND VGND VPWR VPWR U$$853/A sky130_fd_sc_hd__a22o_1
XU$$863 U$$863/A U$$959/A VGND VGND VPWR VPWR U$$863/X sky130_fd_sc_hd__xor2_1
XU$$1002 U$$1002/A U$$992/B VGND VGND VPWR VPWR U$$1002/X sky130_fd_sc_hd__xor2_1
XU$$874 U$$50/B1 U$$910/A2 U$$876/A1 U$$910/B2 VGND VGND VPWR VPWR U$$875/A sky130_fd_sc_hd__a22o_1
XU$$1013 U$$876/A1 U$$999/A2 U$$878/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1014/A sky130_fd_sc_hd__a22o_1
XU$$885 U$$885/A U$$923/B VGND VGND VPWR VPWR U$$885/X sky130_fd_sc_hd__xor2_1
XU$$1024 U$$1024/A U$$980/B VGND VGND VPWR VPWR U$$1024/X sky130_fd_sc_hd__xor2_1
XFILLER_90_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1035 U$$76/A1 U$$1093/A2 U$$76/B1 U$$1073/B2 VGND VGND VPWR VPWR U$$1036/A sky130_fd_sc_hd__a22o_1
XU$$896 U$$74/A1 U$$910/A2 U$$76/A1 U$$910/B2 VGND VGND VPWR VPWR U$$897/A sky130_fd_sc_hd__a22o_1
X_722__774 VGND VGND VPWR VPWR _722__774/HI U$$1650/A1 sky130_fd_sc_hd__conb_1
XU$$1046 U$$1046/A U$$980/B VGND VGND VPWR VPWR U$$1046/X sky130_fd_sc_hd__xor2_1
XU$$1057 U$$96/B1 U$$1093/A2 U$$785/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1058/A sky130_fd_sc_hd__a22o_1
XFILLER_189_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1068 U$$1068/A U$$998/B VGND VGND VPWR VPWR U$$1068/X sky130_fd_sc_hd__xor2_1
XFILLER_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1079 U$$942/A1 U$$963/X U$$944/A1 U$$964/X VGND VGND VPWR VPWR U$$1080/A sky130_fd_sc_hd__a22o_1
XFILLER_176_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_98_4 U$$3927/X U$$4060/X U$$4193/X VGND VGND VPWR VPWR dadda_fa_3_99_2/A
+ dadda_fa_3_98_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_41_0 U$$1552/X U$$1685/X U$$1818/X VGND VGND VPWR VPWR dadda_fa_3_42_0/B
+ dadda_fa_3_41_2/B sky130_fd_sc_hd__fa_2
XFILLER_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2270 U$$76/B1 U$$2270/A2 U$$902/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2271/A sky130_fd_sc_hd__a22o_1
XFILLER_179_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2281 U$$2281/A U$$2289/B VGND VGND VPWR VPWR U$$2281/X sky130_fd_sc_hd__xor2_1
XFILLER_168_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2292 U$$4484/A1 U$$2316/A2 _599_/Q U$$2316/B2 VGND VGND VPWR VPWR U$$2293/A sky130_fd_sc_hd__a22o_1
XU$$1580 U$$1580/A U$$1580/B VGND VGND VPWR VPWR U$$1580/X sky130_fd_sc_hd__xor2_1
XFILLER_179_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1591 U$$84/A1 U$$1591/A2 U$$86/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1592/A sky130_fd_sc_hd__a22o_1
XFILLER_148_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_70_2 dadda_fa_4_70_2/A dadda_fa_4_70_2/B dadda_fa_4_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/CIN dadda_fa_5_70_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_2 U$$2307/X U$$2440/X U$$2573/X VGND VGND VPWR VPWR dadda_fa_2_87_3/B
+ dadda_fa_2_86_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_63_1 dadda_fa_4_63_1/A dadda_fa_4_63_1/B dadda_fa_4_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/B dadda_fa_5_63_1/B sky130_fd_sc_hd__fa_1
XFILLER_89_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_79_1 U$$1495/X U$$1628/X U$$1761/X VGND VGND VPWR VPWR dadda_fa_2_80_0/CIN
+ dadda_fa_2_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_40_0 dadda_fa_7_40_0/A dadda_fa_7_40_0/B dadda_fa_7_40_0/CIN VGND VGND
+ VPWR VPWR _465_/D _336_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_56_0 dadda_fa_4_56_0/A dadda_fa_4_56_0/B dadda_fa_4_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/A dadda_fa_5_56_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$210 final_adder.U$$705/A final_adder.U$$704/A VGND VGND VPWR VPWR
+ final_adder.U$$296/A sky130_fd_sc_hd__and2_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$221 final_adder.U$$715/A final_adder.U$$587/B1 final_adder.U$$221/B1
+ VGND VGND VPWR VPWR final_adder.U$$221/X sky130_fd_sc_hd__a21o_1
XFILLER_85_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$232 final_adder.U$$727/A final_adder.U$$726/A VGND VGND VPWR VPWR
+ final_adder.U$$308/B sky130_fd_sc_hd__and2_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$243 final_adder.U$$737/A final_adder.U$$609/B1 final_adder.U$$243/B1
+ VGND VGND VPWR VPWR final_adder.U$$243/X sky130_fd_sc_hd__a21o_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$265 final_adder.U$$264/A final_adder.U$$145/X final_adder.U$$147/X
+ VGND VGND VPWR VPWR final_adder.U$$265/X sky130_fd_sc_hd__a21o_1
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$104 U$$926/A1 U$$4/X U$$928/A1 U$$5/X VGND VGND VPWR VPWR U$$105/A sky130_fd_sc_hd__a22o_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$276 final_adder.U$$276/A final_adder.U$$276/B VGND VGND VPWR VPWR
+ final_adder.U$$330/B sky130_fd_sc_hd__and2_1
X_530_ _532_/CLK _530_/D VGND VGND VPWR VPWR _530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$115 U$$115/A _617_/Q VGND VGND VPWR VPWR U$$115/X sky130_fd_sc_hd__xor2_2
Xrepeater480 U$$2882/X VGND VGND VPWR VPWR U$$2975/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$287 final_adder.U$$286/A final_adder.U$$189/X final_adder.U$$191/X
+ VGND VGND VPWR VPWR final_adder.U$$287/X sky130_fd_sc_hd__a21o_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$126 U$$948/A1 U$$4/X U$$950/A1 U$$5/X VGND VGND VPWR VPWR U$$127/A sky130_fd_sc_hd__a22o_1
Xrepeater491 U$$2316/B2 VGND VGND VPWR VPWR U$$2286/B2 sky130_fd_sc_hd__buf_12
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$298 final_adder.U$$298/A final_adder.U$$298/B VGND VGND VPWR VPWR
+ final_adder.U$$340/A sky130_fd_sc_hd__and2_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$137 U$$89/B VGND VGND VPWR VPWR U$$137/Y sky130_fd_sc_hd__inv_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$148 U$$148/A U$$242/B VGND VGND VPWR VPWR U$$148/X sky130_fd_sc_hd__xor2_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$159 U$$22/A1 U$$141/X _560_/Q U$$142/X VGND VGND VPWR VPWR U$$160/A sky130_fd_sc_hd__a22o_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_461_ _461_/CLK _461_/D VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_392_ _583_/CLK _392_/D VGND VGND VPWR VPWR _392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_74_0 _683__903/HI U$$820/X U$$953/X VGND VGND VPWR VPWR dadda_fa_1_75_7/CIN
+ dadda_fa_1_74_8/B sky130_fd_sc_hd__fa_2
XFILLER_110_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput250 c[94] VGND VGND VPWR VPWR input250/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$660 U$$934/A1 U$$682/A2 U$$799/A1 U$$553/X VGND VGND VPWR VPWR U$$661/A sky130_fd_sc_hd__a22o_1
X_659_ _667_/CLK _659_/D VGND VGND VPWR VPWR _659_/Q sky130_fd_sc_hd__dfxtp_4
XU$$671 U$$671/A _625_/Q VGND VGND VPWR VPWR U$$671/X sky130_fd_sc_hd__xor2_1
XU$$682 U$$956/A1 U$$682/A2 U$$682/B1 U$$553/X VGND VGND VPWR VPWR U$$683/A sky130_fd_sc_hd__a22o_1
XFILLER_17_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$693 _552_/Q U$$689/X U$$969/A1 U$$817/B2 VGND VGND VPWR VPWR U$$694/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_80_1 dadda_fa_5_80_1/A dadda_fa_5_80_1/B dadda_fa_5_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/B dadda_fa_7_80_0/A sky130_fd_sc_hd__fa_1
XFILLER_160_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_96_1 U$$2859/X U$$2992/X U$$3125/X VGND VGND VPWR VPWR dadda_fa_3_97_0/CIN
+ dadda_fa_3_96_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_73_0 dadda_fa_5_73_0/A dadda_fa_5_73_0/B dadda_fa_5_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/A dadda_fa_6_73_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_89_0 U$$3377/X U$$3510/X U$$3643/X VGND VGND VPWR VPWR dadda_fa_3_90_0/B
+ dadda_fa_3_89_2/B sky130_fd_sc_hd__fa_2
XFILLER_63_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_72_8 dadda_fa_1_72_8/A dadda_fa_1_72_8/B dadda_fa_1_72_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_3/A dadda_fa_3_72_0/A sky130_fd_sc_hd__fa_2
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_65_7 dadda_fa_1_65_7/A dadda_fa_1_65_7/B dadda_fa_1_65_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/CIN dadda_fa_2_65_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_6 U$$3980/X U$$4044/B input210/X VGND VGND VPWR VPWR dadda_fa_2_59_2/B
+ dadda_fa_2_58_5/B sky130_fd_sc_hd__fa_2
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_92_2 U$$2718/X U$$2851/X VGND VGND VPWR VPWR dadda_fa_2_93_5/B dadda_fa_3_92_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_167_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_88_0 dadda_fa_7_88_0/A dadda_fa_7_88_0/B dadda_fa_7_88_0/CIN VGND VGND
+ VPWR VPWR _513_/D _384_/D sky130_fd_sc_hd__fa_1
XFILLER_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_91_0 U$$1917/Y U$$2051/X U$$2184/X VGND VGND VPWR VPWR dadda_fa_2_92_4/B
+ dadda_fa_2_91_5/B sky130_fd_sc_hd__fa_2
XFILLER_117_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4408 _560_/Q U$$4388/X _561_/Q U$$4389/X VGND VGND VPWR VPWR U$$4409/A sky130_fd_sc_hd__a22o_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4419 U$$4419/A U$$4419/B VGND VGND VPWR VPWR U$$4419/X sky130_fd_sc_hd__xor2_2
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3707 U$$4255/A1 U$$3783/A2 U$$969/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3708/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3718 U$$3718/A U$$3756/B VGND VGND VPWR VPWR U$$3718/X sky130_fd_sc_hd__xor2_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3729 _563_/Q U$$3783/A2 _564_/Q U$$3783/B2 VGND VGND VPWR VPWR U$$3730/A sky130_fd_sc_hd__a22o_1
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_103_0 dadda_fa_6_103_0/A dadda_fa_6_103_0/B dadda_fa_6_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_104_0/B dadda_fa_7_103_0/CIN sky130_fd_sc_hd__fa_2
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ _518_/CLK _513_/D VGND VGND VPWR VPWR _513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_23_3 U$$1516/X input172/X dadda_fa_3_23_3/CIN VGND VGND VPWR VPWR dadda_fa_4_24_1/B
+ dadda_fa_4_23_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_444_ _452_/CLK _444_/D VGND VGND VPWR VPWR _444_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_375_ _509_/CLK _375_/D VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_793__845 VGND VGND VPWR VPWR _793__845/HI U$$4431/B sky130_fd_sc_hd__conb_1
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_90_0 dadda_fa_6_90_0/A dadda_fa_6_90_0/B dadda_fa_6_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_91_0/B dadda_fa_7_90_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_834__886 VGND VGND VPWR VPWR _834__886/HI U$$4513/B sky130_fd_sc_hd__conb_1
XFILLER_103_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_5 dadda_fa_2_68_5/A dadda_fa_2_68_5/B dadda_fa_2_68_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_2/A dadda_fa_4_68_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_728__780 VGND VGND VPWR VPWR _728__780/HI U$$2061/A1 sky130_fd_sc_hd__conb_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$490 U$$490/A U$$530/B VGND VGND VPWR VPWR U$$490/X sky130_fd_sc_hd__xor2_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_70_5 U$$4270/X U$$4403/X input224/X VGND VGND VPWR VPWR dadda_fa_2_71_2/A
+ dadda_fa_2_70_5/A sky130_fd_sc_hd__fa_2
XFILLER_8_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_4 U$$3990/X U$$4123/X U$$4256/X VGND VGND VPWR VPWR dadda_fa_2_64_1/CIN
+ dadda_fa_2_63_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_56_3 U$$2380/X U$$2513/X U$$2646/X VGND VGND VPWR VPWR dadda_fa_2_57_1/B
+ dadda_fa_2_56_4/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_33_2 dadda_fa_4_33_2/A dadda_fa_4_33_2/B dadda_fa_4_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/CIN dadda_fa_5_33_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_2 U$$903/X U$$1036/X U$$1169/X VGND VGND VPWR VPWR dadda_fa_2_50_1/B
+ dadda_fa_2_49_4/B sky130_fd_sc_hd__fa_1
XFILLER_43_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_26_1 dadda_fa_4_26_1/A dadda_fa_4_26_1/B dadda_fa_4_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/B dadda_fa_5_26_1/B sky130_fd_sc_hd__fa_1
XFILLER_131_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_0 U$$1109/X U$$1242/X input167/X VGND VGND VPWR VPWR dadda_fa_5_20_0/A
+ dadda_fa_5_19_1/A sky130_fd_sc_hd__fa_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_777__829 VGND VGND VPWR VPWR _777__829/HI U$$4399/B sky130_fd_sc_hd__conb_1
XFILLER_39_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4205 U$$4205/A _677_/Q VGND VGND VPWR VPWR U$$4205/X sky130_fd_sc_hd__xor2_1
XFILLER_77_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4216 U$$654/A1 U$$4244/A2 U$$4492/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4217/A
+ sky130_fd_sc_hd__a22o_1
XU$$4227 U$$4227/A U$$4246/A VGND VGND VPWR VPWR U$$4227/X sky130_fd_sc_hd__xor2_1
XFILLER_59_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4238 U$$539/A1 U$$4244/A2 _613_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4239/A sky130_fd_sc_hd__a22o_1
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3504 U$$3504/A _667_/Q VGND VGND VPWR VPWR U$$3504/X sky130_fd_sc_hd__xor2_1
XU$$4249 U$$4332/B VGND VGND VPWR VPWR U$$4249/Y sky130_fd_sc_hd__inv_1
XU$$3515 _593_/Q U$$3545/A2 _594_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3516/A sky130_fd_sc_hd__a22o_1
XFILLER_19_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3526 U$$3526/A U$$3536/B VGND VGND VPWR VPWR U$$3526/X sky130_fd_sc_hd__xor2_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3537 U$$4496/A1 U$$3429/X U$$936/A1 U$$3430/X VGND VGND VPWR VPWR U$$3538/A sky130_fd_sc_hd__a22o_1
XU$$3548 U$$3548/A U$$3561/A VGND VGND VPWR VPWR U$$3548/X sky130_fd_sc_hd__xor2_1
XU$$2803 U$$2803/A U$$2839/B VGND VGND VPWR VPWR U$$2803/X sky130_fd_sc_hd__xor2_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2814 _585_/Q U$$2870/A2 _586_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2815/A sky130_fd_sc_hd__a22o_1
XU$$3559 U$$819/A1 U$$3429/X U$$3559/B1 U$$3430/X VGND VGND VPWR VPWR U$$3560/A sky130_fd_sc_hd__a22o_1
XFILLER_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2825 U$$2825/A U$$2839/B VGND VGND VPWR VPWR U$$2825/X sky130_fd_sc_hd__xor2_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2836 U$$94/B1 U$$2868/A2 _597_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2837/A sky130_fd_sc_hd__a22o_1
XFILLER_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_21_0 U$$49/X U$$182/X U$$315/X VGND VGND VPWR VPWR dadda_fa_4_22_0/B dadda_fa_4_21_1/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_61_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2847 U$$2847/A U$$2871/B VGND VGND VPWR VPWR U$$2847/X sky130_fd_sc_hd__xor2_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2858 _607_/Q U$$2870/A2 _608_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2859/A sky130_fd_sc_hd__a22o_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2869 U$$2869/A U$$2871/B VGND VGND VPWR VPWR U$$2869/X sky130_fd_sc_hd__xor2_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ _438_/CLK _427_/D VGND VGND VPWR VPWR _427_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_358_ _492_/CLK _358_/D VGND VGND VPWR VPWR _358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_289_ _612_/CLK _289_/D VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_80_4 dadda_fa_2_80_4/A dadda_fa_2_80_4/B dadda_fa_2_80_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/CIN dadda_fa_3_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_73_3 dadda_fa_2_73_3/A dadda_fa_2_73_3/B dadda_fa_2_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/B dadda_fa_3_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_64_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_66_2 dadda_fa_2_66_2/A dadda_fa_2_66_2/B dadda_fa_2_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/A dadda_fa_3_66_3/A sky130_fd_sc_hd__fa_2
XFILLER_122_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_43_1 dadda_fa_5_43_1/A dadda_fa_5_43_1/B dadda_fa_5_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/B dadda_fa_7_43_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_59_1 dadda_fa_2_59_1/A dadda_fa_2_59_1/B dadda_fa_2_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/CIN dadda_fa_3_59_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 a[11] VGND VGND VPWR VPWR _627_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_49_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_36_0 dadda_fa_5_36_0/A dadda_fa_5_36_0/B dadda_fa_5_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/A dadda_fa_6_36_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_25_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_110_0 dadda_fa_5_110_0/A dadda_fa_5_110_0/B dadda_fa_5_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/A dadda_fa_6_110_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1 _425_/Q _297_/Q VGND VGND VPWR VPWR final_adder.U$$129/B1 final_adder.U$$623/A
+ sky130_fd_sc_hd__ha_1
XFILLER_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput340 _173_/Q VGND VGND VPWR VPWR o[5] sky130_fd_sc_hd__buf_2
XFILLER_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput351 _174_/Q VGND VGND VPWR VPWR o[6] sky130_fd_sc_hd__buf_2
Xoutput362 _175_/Q VGND VGND VPWR VPWR o[7] sky130_fd_sc_hd__buf_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput373 _176_/Q VGND VGND VPWR VPWR o[8] sky130_fd_sc_hd__buf_2
XFILLER_114_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput384 _177_/Q VGND VGND VPWR VPWR o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_61_1 U$$2390/X U$$2523/X U$$2656/X VGND VGND VPWR VPWR dadda_fa_2_62_0/CIN
+ dadda_fa_2_61_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_54_0 U$$780/X U$$913/X U$$1046/X VGND VGND VPWR VPWR dadda_fa_2_55_0/B
+ dadda_fa_2_54_3/B sky130_fd_sc_hd__fa_1
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1409 U$$1409/A U$$1461/B VGND VGND VPWR VPWR U$$1409/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_212_ _456_/CLK _212_/D VGND VGND VPWR VPWR _212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_90_3 dadda_fa_3_90_3/A dadda_fa_3_90_3/B dadda_fa_3_90_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/B dadda_fa_4_90_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_109_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_83_2 dadda_fa_3_83_2/A dadda_fa_3_83_2/B dadda_fa_3_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/A dadda_fa_4_83_2/B sky130_fd_sc_hd__fa_1
XFILLER_48_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_76_1 dadda_fa_3_76_1/A dadda_fa_3_76_1/B dadda_fa_3_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/CIN dadda_fa_4_76_2/A sky130_fd_sc_hd__fa_1
XFILLER_151_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_53_0 dadda_fa_6_53_0/A dadda_fa_6_53_0/B dadda_fa_6_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_54_0/B dadda_fa_7_53_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_69_0 dadda_fa_3_69_0/A dadda_fa_3_69_0/B dadda_fa_3_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/B dadda_fa_4_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4002 U$$4002/A U$$4058/B VGND VGND VPWR VPWR U$$4002/X sky130_fd_sc_hd__xor2_1
XU$$4013 U$$4424/A1 U$$4107/A2 _569_/Q U$$4107/B2 VGND VGND VPWR VPWR U$$4014/A sky130_fd_sc_hd__a22o_1
XFILLER_93_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4024 U$$4024/A U$$4058/B VGND VGND VPWR VPWR U$$4024/X sky130_fd_sc_hd__xor2_1
XFILLER_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4035 U$$4446/A1 U$$4045/A2 _580_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$4036/A sky130_fd_sc_hd__a22o_1
XFILLER_24_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4046 U$$4046/A _675_/Q VGND VGND VPWR VPWR U$$4046/X sky130_fd_sc_hd__xor2_1
XU$$3301 U$$3301/A U$$3397/B VGND VGND VPWR VPWR U$$3301/X sky130_fd_sc_hd__xor2_1
XU$$3312 _560_/Q U$$3412/A2 _561_/Q U$$3412/B2 VGND VGND VPWR VPWR U$$3313/A sky130_fd_sc_hd__a22o_1
XU$$4057 _590_/Q U$$3977/X U$$908/A1 U$$3978/X VGND VGND VPWR VPWR U$$4058/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_112_2 dadda_fa_4_112_2/A dadda_fa_4_112_2/B dadda_ha_3_112_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/CIN dadda_fa_5_112_1/CIN sky130_fd_sc_hd__fa_1
XU$$4068 U$$4068/A _675_/Q VGND VGND VPWR VPWR U$$4068/X sky130_fd_sc_hd__xor2_1
XU$$3323 U$$3323/A U$$3397/B VGND VGND VPWR VPWR U$$3323/X sky130_fd_sc_hd__xor2_1
XFILLER_81_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3334 U$$4291/B1 U$$3396/A2 U$$4156/B1 U$$3396/B2 VGND VGND VPWR VPWR U$$3335/A
+ sky130_fd_sc_hd__a22o_1
XU$$4079 U$$654/A1 U$$4107/A2 U$$4492/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4080/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3345 U$$3345/A U$$3403/B VGND VGND VPWR VPWR U$$3345/X sky130_fd_sc_hd__xor2_1
XU$$2600 U$$956/A1 U$$2470/X U$$2600/B1 U$$2471/X VGND VGND VPWR VPWR U$$2601/A sky130_fd_sc_hd__a22o_1
XU$$2611 U$$8/A1 U$$2729/A2 U$$8/B1 U$$2729/B2 VGND VGND VPWR VPWR U$$2612/A sky130_fd_sc_hd__a22o_1
XU$$3356 _582_/Q U$$3412/A2 U$$70/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3357/A sky130_fd_sc_hd__a22o_1
XU$$3367 U$$3367/A U$$3403/B VGND VGND VPWR VPWR U$$3367/X sky130_fd_sc_hd__xor2_1
XU$$2622 U$$2622/A U$$2694/B VGND VGND VPWR VPWR U$$2622/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_105_1 dadda_fa_4_105_1/A dadda_fa_4_105_1/B dadda_fa_4_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/B dadda_fa_5_105_1/B sky130_fd_sc_hd__fa_1
XFILLER_74_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3378 _593_/Q U$$3292/X _594_/Q U$$3293/X VGND VGND VPWR VPWR U$$3379/A sky130_fd_sc_hd__a22o_1
XU$$2633 U$$30/A1 U$$2667/A2 U$$30/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2634/A sky130_fd_sc_hd__a22o_1
XFILLER_19_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2644 U$$2644/A U$$2694/B VGND VGND VPWR VPWR U$$2644/X sky130_fd_sc_hd__xor2_1
X_799__851 VGND VGND VPWR VPWR _799__851/HI U$$4443/B sky130_fd_sc_hd__conb_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1910 U$$1910/A _643_/Q VGND VGND VPWR VPWR U$$1910/X sky130_fd_sc_hd__xor2_1
XU$$3389 U$$3389/A U$$3403/B VGND VGND VPWR VPWR U$$3389/X sky130_fd_sc_hd__xor2_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2655 U$$2790/B1 U$$2667/A2 U$$876/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2656/A
+ sky130_fd_sc_hd__a22o_1
XU$$1921 U$$2055/A U$$1921/B VGND VGND VPWR VPWR U$$1921/X sky130_fd_sc_hd__and2_1
XU$$2666 U$$2666/A U$$2710/B VGND VGND VPWR VPWR U$$2666/X sky130_fd_sc_hd__xor2_1
XU$$2677 U$$4045/B1 U$$2607/X _586_/Q U$$2608/X VGND VGND VPWR VPWR U$$2678/A sky130_fd_sc_hd__a22o_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1932 U$$14/A1 U$$2048/A2 U$$14/B1 U$$2048/B2 VGND VGND VPWR VPWR U$$1933/A sky130_fd_sc_hd__a22o_1
XU$$2688 U$$2688/A U$$2698/B VGND VGND VPWR VPWR U$$2688/X sky130_fd_sc_hd__xor2_1
XU$$1943 U$$1943/A U$$2021/B VGND VGND VPWR VPWR U$$1943/X sky130_fd_sc_hd__xor2_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2699 _596_/Q U$$2607/X _597_/Q U$$2608/X VGND VGND VPWR VPWR U$$2700/A sky130_fd_sc_hd__a22o_1
XU$$1954 U$$4283/A1 U$$2036/A2 U$$4285/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1955/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1965 U$$1965/A U$$2023/B VGND VGND VPWR VPWR U$$1965/X sky130_fd_sc_hd__xor2_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1976 U$$880/A1 U$$2036/A2 U$$4170/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1977/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1987 U$$1987/A U$$2023/B VGND VGND VPWR VPWR U$$1987/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_126_0 dadda_fa_7_126_0/A dadda_fa_7_126_0/B dadda_fa_7_126_0/CIN VGND
+ VGND VPWR VPWR _551_/D _422_/D sky130_fd_sc_hd__fa_1
XU$$1998 U$$765/A1 U$$2052/A2 U$$82/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$1999/A sky130_fd_sc_hd__a22o_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_71_0 dadda_fa_2_71_0/A dadda_fa_2_71_0/B dadda_fa_2_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/B dadda_fa_3_71_2/B sky130_fd_sc_hd__fa_2
XFILLER_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$617 final_adder.U$$744/A final_adder.U$$744/B final_adder.U$$617/B1
+ VGND VGND VPWR VPWR final_adder.U$$745/B sky130_fd_sc_hd__a21o_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$628 final_adder.U$$628/A final_adder.U$$628/B VGND VGND VPWR VPWR
+ _174_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$639 final_adder.U$$639/A final_adder.U$$639/B VGND VGND VPWR VPWR
+ _185_/D sky130_fd_sc_hd__xor2_1
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$50 U$$50/A1 U$$4/X U$$50/B1 U$$5/X VGND VGND VPWR VPWR U$$51/A sky130_fd_sc_hd__a22o_1
XU$$61 U$$61/A U$$3/A VGND VGND VPWR VPWR U$$61/X sky130_fd_sc_hd__xor2_2
XFILLER_38_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$72 U$$72/A1 U$$4/X U$$74/A1 U$$5/X VGND VGND VPWR VPWR U$$73/A sky130_fd_sc_hd__a22o_1
XU$$83 U$$83/A U$$89/B VGND VGND VPWR VPWR U$$83/X sky130_fd_sc_hd__xor2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$94 U$$94/A1 U$$4/X U$$94/B1 U$$5/X VGND VGND VPWR VPWR U$$95/A sky130_fd_sc_hd__a22o_1
XU$$3890 U$$4438/A1 U$$3840/X U$$4303/A1 U$$3841/X VGND VGND VPWR VPWR U$$3891/A sky130_fd_sc_hd__a22o_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_93_1 dadda_fa_4_93_1/A dadda_fa_4_93_1/B dadda_fa_4_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/B dadda_fa_5_93_1/B sky130_fd_sc_hd__fa_1
XFILLER_137_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_70_0 dadda_fa_7_70_0/A dadda_fa_7_70_0/B dadda_fa_7_70_0/CIN VGND VGND
+ VPWR VPWR _495_/D _366_/D sky130_fd_sc_hd__fa_2
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_86_0 dadda_fa_4_86_0/A dadda_fa_4_86_0/B dadda_fa_4_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/A dadda_fa_5_86_1/A sky130_fd_sc_hd__fa_1
XFILLER_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_107_3 input137/X dadda_fa_3_107_3/B dadda_fa_3_107_3/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_108_1/B dadda_fa_4_107_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1206 _603_/Q U$$1218/A2 _604_/Q U$$1218/B2 VGND VGND VPWR VPWR U$$1207/A sky130_fd_sc_hd__a22o_1
XFILLER_16_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1217 U$$1217/A _633_/Q VGND VGND VPWR VPWR U$$1217/X sky130_fd_sc_hd__xor2_1
XU$$1228 U$$952/B1 U$$1100/X U$$819/A1 U$$1101/X VGND VGND VPWR VPWR U$$1229/A sky130_fd_sc_hd__a22o_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1239 U$$1239/A1 U$$1237/X _552_/Q U$$1238/X VGND VGND VPWR VPWR U$$1240/A sky130_fd_sc_hd__a22o_1
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_50_5 dadda_fa_2_50_5/A dadda_fa_2_50_5/B dadda_fa_2_50_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_2/A dadda_fa_4_50_0/A sky130_fd_sc_hd__fa_2
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_43_4 dadda_fa_2_43_4/A dadda_fa_2_43_4/B dadda_fa_2_43_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/CIN dadda_fa_3_43_3/CIN sky130_fd_sc_hd__fa_1
XU$$3120 U$$654/A1 U$$3146/A2 U$$930/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3121/A sky130_fd_sc_hd__a22o_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3131 U$$3131/A U$$3137/B VGND VGND VPWR VPWR U$$3131/X sky130_fd_sc_hd__xor2_1
XU$$3142 U$$950/A1 U$$3146/A2 U$$4514/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3143/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_6_2_0 U$$11/X U$$144/X VGND VGND VPWR VPWR dadda_fa_7_3_0/B dadda_ha_6_2_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3153 _663_/Q VGND VGND VPWR VPWR U$$3153/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_3 U$$1941/X U$$2074/X U$$2207/X VGND VGND VPWR VPWR dadda_fa_3_37_1/B
+ dadda_fa_3_36_3/B sky130_fd_sc_hd__fa_2
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3164 U$$3164/A U$$3224/B VGND VGND VPWR VPWR U$$3164/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3175 _560_/Q U$$3241/A2 _561_/Q U$$3253/B2 VGND VGND VPWR VPWR U$$3176/A sky130_fd_sc_hd__a22o_1
XU$$2430 U$$2430/A _651_/Q VGND VGND VPWR VPWR U$$2430/X sky130_fd_sc_hd__xor2_1
XU$$2441 U$$934/A1 U$$2463/A2 U$$936/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2442/A sky130_fd_sc_hd__a22o_1
XU$$3186 U$$3186/A U$$3224/B VGND VGND VPWR VPWR U$$3186/X sky130_fd_sc_hd__xor2_2
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3197 U$$46/A1 U$$3241/A2 _572_/Q U$$3253/B2 VGND VGND VPWR VPWR U$$3198/A sky130_fd_sc_hd__a22o_1
XU$$2452 U$$2452/A _651_/Q VGND VGND VPWR VPWR U$$2452/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_29_2 U$$863/X U$$996/X U$$1129/X VGND VGND VPWR VPWR dadda_fa_3_30_2/A
+ dadda_fa_3_29_3/CIN sky130_fd_sc_hd__fa_1
XU$$2463 U$$956/A1 U$$2463/A2 U$$2463/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2464/A
+ sky130_fd_sc_hd__a22o_1
XU$$2474 U$$8/A1 U$$2574/A2 U$$969/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2475/A sky130_fd_sc_hd__a22o_1
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1740 U$$94/B1 U$$1648/X U$$98/A1 U$$1649/X VGND VGND VPWR VPWR U$$1741/A sky130_fd_sc_hd__a22o_1
XU$$2485 U$$2485/A U$$2533/B VGND VGND VPWR VPWR U$$2485/X sky130_fd_sc_hd__xor2_1
XU$$1751 U$$1751/A _641_/Q VGND VGND VPWR VPWR U$$1751/X sky130_fd_sc_hd__xor2_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2496 U$$30/A1 U$$2574/A2 U$$30/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2497/A sky130_fd_sc_hd__a22o_1
XU$$1762 U$$940/A1 U$$1648/X U$$4504/A1 U$$1649/X VGND VGND VPWR VPWR U$$1763/A sky130_fd_sc_hd__a22o_1
XU$$1773 U$$1773/A U$$1781/A VGND VGND VPWR VPWR U$$1773/X sky130_fd_sc_hd__xor2_1
XU$$1784 U$$1918/A U$$1784/B VGND VGND VPWR VPWR U$$1784/X sky130_fd_sc_hd__and2_1
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1795 U$$12/B1 U$$1867/A2 U$$16/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1796/A sky130_fd_sc_hd__a22o_1
XFILLER_148_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput50 a[54] VGND VGND VPWR VPWR _670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput61 a[6] VGND VGND VPWR VPWR _622_/D sky130_fd_sc_hd__buf_4
Xinput72 b[16] VGND VGND VPWR VPWR _568_/D sky130_fd_sc_hd__buf_2
Xinput83 b[26] VGND VGND VPWR VPWR _578_/D sky130_fd_sc_hd__buf_2
Xinput94 b[36] VGND VGND VPWR VPWR _588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$403 final_adder.U$$348/X final_adder.U$$734/B final_adder.U$$349/X
+ VGND VGND VPWR VPWR final_adder.U$$742/B sky130_fd_sc_hd__a21o_2
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$425 final_adder.U$$342/B final_adder.U$$710/B final_adder.U$$301/X
+ VGND VGND VPWR VPWR final_adder.U$$714/B sky130_fd_sc_hd__a21o_1
XFILLER_123_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater640 _602_/Q VGND VGND VPWR VPWR U$$928/B1 sky130_fd_sc_hd__buf_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$447 final_adder.U$$270/B final_adder.U$$650/B final_adder.U$$157/X
+ VGND VGND VPWR VPWR final_adder.U$$652/B sky130_fd_sc_hd__a21o_1
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater651 _597_/Q VGND VGND VPWR VPWR U$$96/B1 sky130_fd_sc_hd__buf_12
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater662 U$$4335/A1 VGND VGND VPWR VPWR U$$771/B1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$469 final_adder.U$$292/B final_adder.U$$694/B final_adder.U$$201/X
+ VGND VGND VPWR VPWR final_adder.U$$696/B sky130_fd_sc_hd__a21o_1
XU$$308 U$$34/A1 U$$278/X U$$36/A1 U$$279/X VGND VGND VPWR VPWR U$$309/A sky130_fd_sc_hd__a22o_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater673 U$$765/A1 VGND VGND VPWR VPWR U$$80/A1 sky130_fd_sc_hd__buf_12
XFILLER_26_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$319 U$$319/A U$$357/B VGND VGND VPWR VPWR U$$319/X sky130_fd_sc_hd__xor2_1
Xrepeater684 _584_/Q VGND VGND VPWR VPWR U$$892/B1 sky130_fd_sc_hd__buf_12
Xrepeater695 _580_/Q VGND VGND VPWR VPWR U$$3900/A1 sky130_fd_sc_hd__buf_12
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_112_1 U$$3689/X U$$3822/X U$$3955/X VGND VGND VPWR VPWR dadda_fa_4_113_1/CIN
+ dadda_fa_4_112_2/B sky130_fd_sc_hd__fa_1
XFILLER_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_105_0 U$$3675/X U$$3808/X U$$3941/X VGND VGND VPWR VPWR dadda_fa_4_106_0/B
+ dadda_fa_4_105_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_53_3 dadda_fa_3_53_3/A dadda_fa_3_53_3/B dadda_fa_3_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/B dadda_fa_4_53_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_69_3 U$$1608/X U$$1741/X U$$1874/X VGND VGND VPWR VPWR dadda_fa_1_70_7/A
+ dadda_fa_1_69_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_46_2 dadda_fa_3_46_2/A dadda_fa_3_46_2/B dadda_fa_3_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/A dadda_fa_4_46_2/B sky130_fd_sc_hd__fa_1
XFILLER_91_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$820 U$$820/A U$$822/A VGND VGND VPWR VPWR U$$820/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_39_1 dadda_fa_3_39_1/A dadda_fa_3_39_1/B dadda_fa_3_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/CIN dadda_fa_4_39_2/A sky130_fd_sc_hd__fa_2
X_675_ _678_/CLK _675_/D VGND VGND VPWR VPWR _675_/Q sky130_fd_sc_hd__dfxtp_4
XU$$831 U$$831/A U$$923/B VGND VGND VPWR VPWR U$$831/X sky130_fd_sc_hd__xor2_1
XFILLER_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$842 U$$842/A1 U$$928/A2 U$$22/A1 U$$928/B2 VGND VGND VPWR VPWR U$$843/A sky130_fd_sc_hd__a22o_1
XFILLER_189_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_16_0 dadda_fa_6_16_0/A dadda_fa_6_16_0/B dadda_fa_6_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_17_0/B dadda_fa_7_16_0/CIN sky130_fd_sc_hd__fa_1
XU$$853 U$$853/A U$$903/B VGND VGND VPWR VPWR U$$853/X sky130_fd_sc_hd__xor2_1
XU$$1003 U$$4291/A1 U$$999/A2 U$$868/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1004/A sky130_fd_sc_hd__a22o_1
XFILLER_189_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$864 _569_/Q U$$928/A2 _570_/Q U$$928/B2 VGND VGND VPWR VPWR U$$865/A sky130_fd_sc_hd__a22o_1
XU$$875 U$$875/A U$$903/B VGND VGND VPWR VPWR U$$875/X sky130_fd_sc_hd__xor2_1
XU$$1014 U$$1014/A U$$980/B VGND VGND VPWR VPWR U$$1014/X sky130_fd_sc_hd__xor2_1
XFILLER_32_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$886 U$$64/A1 U$$928/A2 U$$66/A1 U$$928/B2 VGND VGND VPWR VPWR U$$887/A sky130_fd_sc_hd__a22o_1
XU$$1025 U$$3489/B1 U$$999/A2 U$$3217/B1 U$$987/B2 VGND VGND VPWR VPWR U$$1026/A sky130_fd_sc_hd__a22o_1
XU$$897 U$$897/A U$$903/B VGND VGND VPWR VPWR U$$897/X sky130_fd_sc_hd__xor2_1
XU$$1036 U$$1036/A U$$980/B VGND VGND VPWR VPWR U$$1036/X sky130_fd_sc_hd__xor2_1
XFILLER_189_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1047 U$$88/A1 U$$1093/A2 U$$912/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1048/A sky130_fd_sc_hd__a22o_1
XFILLER_189_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1058 U$$1058/A U$$980/B VGND VGND VPWR VPWR U$$1058/X sky130_fd_sc_hd__xor2_1
XU$$1069 U$$932/A1 U$$963/X U$$934/A1 U$$964/X VGND VGND VPWR VPWR U$$1070/A sky130_fd_sc_hd__a22o_1
XFILLER_176_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_41_1 U$$1951/X U$$2084/X U$$2217/X VGND VGND VPWR VPWR dadda_fa_3_42_0/CIN
+ dadda_fa_3_41_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_34_0 U$$341/X U$$474/X U$$607/X VGND VGND VPWR VPWR dadda_fa_3_35_0/B
+ dadda_fa_3_34_2/B sky130_fd_sc_hd__fa_2
XFILLER_81_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2260 _582_/Q U$$2196/X U$$70/A1 U$$2197/X VGND VGND VPWR VPWR U$$2261/A sky130_fd_sc_hd__a22o_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2271 U$$2271/A U$$2289/B VGND VGND VPWR VPWR U$$2271/X sky130_fd_sc_hd__xor2_1
XFILLER_168_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2282 _593_/Q U$$2326/A2 _594_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2283/A sky130_fd_sc_hd__a22o_1
XU$$2293 U$$2293/A U$$2327/B VGND VGND VPWR VPWR U$$2293/X sky130_fd_sc_hd__xor2_1
XU$$1570 U$$1570/A U$$1614/B VGND VGND VPWR VPWR U$$1570/X sky130_fd_sc_hd__xor2_1
XU$$1581 U$$74/A1 U$$1605/A2 U$$2953/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1582/A sky130_fd_sc_hd__a22o_1
XFILLER_33_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1592 U$$1592/A U$$1614/B VGND VGND VPWR VPWR U$$1592/X sky130_fd_sc_hd__xor2_1
XFILLER_148_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_86_3 U$$2706/X U$$2839/X U$$2972/X VGND VGND VPWR VPWR dadda_fa_2_87_3/CIN
+ dadda_fa_2_86_5/B sky130_fd_sc_hd__fa_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_63_2 dadda_fa_4_63_2/A dadda_fa_4_63_2/B dadda_fa_4_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/CIN dadda_fa_5_63_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_2 U$$1894/X U$$2027/X U$$2160/X VGND VGND VPWR VPWR dadda_fa_2_80_1/A
+ dadda_fa_2_79_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_56_1 dadda_fa_4_56_1/A dadda_fa_4_56_1/B dadda_fa_4_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/B dadda_fa_5_56_1/B sky130_fd_sc_hd__fa_1
XFILLER_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$200 final_adder.U$$695/A final_adder.U$$694/A VGND VGND VPWR VPWR
+ final_adder.U$$292/B sky130_fd_sc_hd__and2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$211 final_adder.U$$705/A final_adder.U$$577/B1 final_adder.U$$211/B1
+ VGND VGND VPWR VPWR final_adder.U$$211/X sky130_fd_sc_hd__a21o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk _632_/CLK VGND VGND VPWR VPWR _620_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_33_0 dadda_fa_7_33_0/A dadda_fa_7_33_0/B dadda_fa_7_33_0/CIN VGND VGND
+ VPWR VPWR _458_/D _329_/D sky130_fd_sc_hd__fa_2
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$222 final_adder.U$$717/A final_adder.U$$716/A VGND VGND VPWR VPWR
+ final_adder.U$$302/A sky130_fd_sc_hd__and2_1
Xdadda_fa_4_49_0 dadda_fa_4_49_0/A dadda_fa_4_49_0/B dadda_fa_4_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/A dadda_fa_5_49_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$233 final_adder.U$$727/A final_adder.U$$599/B1 final_adder.U$$233/B1
+ VGND VGND VPWR VPWR final_adder.U$$233/X sky130_fd_sc_hd__a21o_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$244 final_adder.U$$739/A final_adder.U$$738/A VGND VGND VPWR VPWR
+ final_adder.U$$314/B sky130_fd_sc_hd__and2_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$266 final_adder.U$$266/A final_adder.U$$266/B VGND VGND VPWR VPWR
+ final_adder.U$$324/A sky130_fd_sc_hd__and2_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$105 U$$105/A U$$3/A VGND VGND VPWR VPWR U$$105/X sky130_fd_sc_hd__xor2_2
Xrepeater470 U$$3668/B2 VGND VGND VPWR VPWR U$$3678/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$277 final_adder.U$$276/A final_adder.U$$169/X final_adder.U$$171/X
+ VGND VGND VPWR VPWR final_adder.U$$277/X sky130_fd_sc_hd__a21o_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$116 U$$938/A1 U$$4/X U$$940/A1 U$$5/X VGND VGND VPWR VPWR U$$117/A sky130_fd_sc_hd__a22o_1
Xrepeater481 U$$2882/X VGND VGND VPWR VPWR U$$3009/B2 sky130_fd_sc_hd__buf_12
XFILLER_84_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$288 final_adder.U$$288/A final_adder.U$$288/B VGND VGND VPWR VPWR
+ final_adder.U$$336/B sky130_fd_sc_hd__and2_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$127 U$$127/A _617_/Q VGND VGND VPWR VPWR U$$127/X sky130_fd_sc_hd__xor2_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater492 U$$2316/B2 VGND VGND VPWR VPWR U$$2326/B2 sky130_fd_sc_hd__buf_12
XFILLER_73_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_745__797 VGND VGND VPWR VPWR _745__797/HI U$$3148/B1 sky130_fd_sc_hd__conb_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$299 final_adder.U$$298/A final_adder.U$$213/X final_adder.U$$215/X
+ VGND VGND VPWR VPWR final_adder.U$$299/X sky130_fd_sc_hd__a21o_1
XU$$138 _618_/Q VGND VGND VPWR VPWR U$$140/B sky130_fd_sc_hd__inv_1
XFILLER_73_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$149 U$$971/A1 U$$141/X U$$12/B1 U$$142/X VGND VGND VPWR VPWR U$$150/A sky130_fd_sc_hd__a22o_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ _462_/CLK _460_/D VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_391_ _535_/CLK _391_/D VGND VGND VPWR VPWR _391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _333_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_74_1 U$$1086/X U$$1219/X U$$1352/X VGND VGND VPWR VPWR dadda_fa_1_75_8/A
+ dadda_fa_1_74_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput240 c[85] VGND VGND VPWR VPWR input240/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_51_0 dadda_fa_3_51_0/A dadda_fa_3_51_0/B dadda_fa_3_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/B dadda_fa_4_51_1/CIN sky130_fd_sc_hd__fa_1
Xinput251 c[95] VGND VGND VPWR VPWR input251/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_67_0 U$$136/Y U$$273/Y U$$407/X VGND VGND VPWR VPWR dadda_fa_1_68_5/B
+ dadda_fa_1_67_7/B sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_87_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _647_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$650 U$$924/A1 U$$682/A2 U$$926/A1 U$$553/X VGND VGND VPWR VPWR U$$651/A sky130_fd_sc_hd__a22o_1
X_658_ _667_/CLK _658_/D VGND VGND VPWR VPWR _658_/Q sky130_fd_sc_hd__dfxtp_1
XU$$661 U$$661/A U$$661/B VGND VGND VPWR VPWR U$$661/X sky130_fd_sc_hd__xor2_1
XFILLER_189_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$672 U$$946/A1 U$$552/X U$$948/A1 U$$553/X VGND VGND VPWR VPWR U$$673/A sky130_fd_sc_hd__a22o_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$683 U$$683/A _625_/Q VGND VGND VPWR VPWR U$$683/X sky130_fd_sc_hd__xor2_1
XU$$694 U$$694/A U$$784/B VGND VGND VPWR VPWR U$$694/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_589_ _597_/CLK _589_/D VGND VGND VPWR VPWR _589_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_694__914 VGND VGND VPWR VPWR _694__914/HI _694__914/LO sky130_fd_sc_hd__conb_1
XFILLER_158_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_11_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _455_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_96_2 U$$3258/X U$$3391/X U$$3524/X VGND VGND VPWR VPWR dadda_fa_3_97_1/A
+ dadda_fa_3_96_3/A sky130_fd_sc_hd__fa_2
XFILLER_133_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_73_1 dadda_fa_5_73_1/A dadda_fa_5_73_1/B dadda_fa_5_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/B dadda_fa_7_73_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_89_1 U$$3776/X U$$3909/X U$$4042/X VGND VGND VPWR VPWR dadda_fa_3_90_0/CIN
+ dadda_fa_3_89_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_125_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_66_0 dadda_fa_5_66_0/A dadda_fa_5_66_0/B dadda_fa_5_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/A dadda_fa_6_66_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_65_8 dadda_fa_1_65_8/A dadda_fa_1_65_8/B dadda_fa_1_65_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_3/A dadda_fa_3_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_78_clk _560_/CLK VGND VGND VPWR VPWR _551_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_7 dadda_fa_1_58_7/A dadda_fa_1_58_7/B dadda_fa_1_58_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_2/CIN dadda_fa_2_58_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_5_0 U$$283/X input212/X dadda_fa_6_5_0/CIN VGND VGND VPWR VPWR dadda_fa_7_6_0/B
+ dadda_fa_7_5_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2090 U$$2090/A U$$2118/B VGND VGND VPWR VPWR U$$2090/X sky130_fd_sc_hd__xor2_1
XFILLER_161_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_91_1 U$$2317/X U$$2450/X U$$2583/X VGND VGND VPWR VPWR dadda_fa_2_92_4/CIN
+ dadda_fa_2_91_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_84_0 _687__907/HI U$$1505/X U$$1638/X VGND VGND VPWR VPWR dadda_fa_2_85_2/A
+ dadda_fa_2_84_4/A sky130_fd_sc_hd__fa_1
XFILLER_2_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4409 U$$4409/A U$$4409/B VGND VGND VPWR VPWR U$$4409/X sky130_fd_sc_hd__xor2_1
XFILLER_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_clk _560_/CLK VGND VGND VPWR VPWR _677_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3708 U$$3708/A U$$3784/B VGND VGND VPWR VPWR U$$3708/X sky130_fd_sc_hd__xor2_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3719 U$$979/A1 U$$3795/A2 U$$22/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3720/A sky130_fd_sc_hd__a22o_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _518_/CLK _512_/D VGND VGND VPWR VPWR _512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _455_/CLK _443_/D VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _503_/CLK _374_/D VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_83_0 dadda_fa_6_83_0/A dadda_fa_6_83_0/B dadda_fa_6_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_84_0/B dadda_fa_7_83_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_99_0 U$$4461/X input255/X dadda_fa_3_99_0/CIN VGND VGND VPWR VPWR dadda_fa_4_100_0/B
+ dadda_fa_4_99_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_0_clk _632_/CLK VGND VGND VPWR VPWR _303_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$480 U$$480/A U$$547/A VGND VGND VPWR VPWR U$$480/X sky130_fd_sc_hd__xor2_1
XU$$491 U$$902/A1 U$$491/A2 U$$902/B1 U$$416/X VGND VGND VPWR VPWR U$$492/A sky130_fd_sc_hd__a22o_1
XFILLER_149_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_70_6 dadda_fa_1_70_6/A dadda_fa_1_70_6/B dadda_fa_1_70_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/B dadda_fa_2_70_5/B sky130_fd_sc_hd__fa_1
XFILLER_113_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_63_5 input216/X dadda_fa_1_63_5/B dadda_fa_1_63_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_64_2/A dadda_fa_2_63_5/A sky130_fd_sc_hd__fa_2
XFILLER_41_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_56_4 U$$2779/X U$$2912/X U$$3045/X VGND VGND VPWR VPWR dadda_fa_2_57_1/CIN
+ dadda_fa_2_56_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_49_3 U$$1302/X U$$1435/X U$$1568/X VGND VGND VPWR VPWR dadda_fa_2_50_1/CIN
+ dadda_fa_2_49_4/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_26_2 dadda_fa_4_26_2/A dadda_fa_4_26_2/B dadda_fa_4_26_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/CIN dadda_fa_5_26_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_1 dadda_fa_4_19_1/A dadda_fa_4_19_1/B dadda_fa_4_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/B dadda_fa_5_19_1/B sky130_fd_sc_hd__fa_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4206 _596_/Q U$$4114/X U$$98/A1 U$$4115/X VGND VGND VPWR VPWR U$$4207/A sky130_fd_sc_hd__a22o_1
XFILLER_59_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4217 U$$4217/A U$$4246/A VGND VGND VPWR VPWR U$$4217/X sky130_fd_sc_hd__xor2_1
XFILLER_93_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4228 U$$4502/A1 U$$4244/A2 U$$4504/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4229/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4239 U$$4239/A U$$4246/A VGND VGND VPWR VPWR U$$4239/X sky130_fd_sc_hd__xor2_1
XU$$3505 U$$765/A1 U$$3545/A2 U$$630/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3506/A sky130_fd_sc_hd__a22o_1
XU$$3516 U$$3516/A U$$3536/B VGND VGND VPWR VPWR U$$3516/X sky130_fd_sc_hd__xor2_1
XFILLER_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3527 U$$4486/A1 U$$3545/A2 U$$787/B1 U$$3545/B2 VGND VGND VPWR VPWR U$$3528/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_760__812 VGND VGND VPWR VPWR _760__812/HI U$$408/B1 sky130_fd_sc_hd__conb_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3538 U$$3538/A U$$3561/A VGND VGND VPWR VPWR U$$3538/X sky130_fd_sc_hd__xor2_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3549 U$$4508/A1 U$$3429/X U$$4510/A1 U$$3430/X VGND VGND VPWR VPWR U$$3550/A sky130_fd_sc_hd__a22o_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2804 U$$3900/A1 U$$2868/A2 U$$3489/B1 U$$2826/B2 VGND VGND VPWR VPWR U$$2805/A
+ sky130_fd_sc_hd__a22o_1
XU$$2815 U$$2815/A U$$2871/B VGND VGND VPWR VPWR U$$2815/X sky130_fd_sc_hd__xor2_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2826 U$$86/A1 U$$2868/A2 U$$88/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2827/A sky130_fd_sc_hd__a22o_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2837 U$$2837/A U$$2871/B VGND VGND VPWR VPWR U$$2837/X sky130_fd_sc_hd__xor2_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2848 U$$928/B1 U$$2870/A2 U$$4494/A1 U$$2870/B2 VGND VGND VPWR VPWR U$$2849/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_1 U$$448/X U$$581/X U$$714/X VGND VGND VPWR VPWR dadda_fa_4_22_0/CIN
+ dadda_fa_4_21_2/A sky130_fd_sc_hd__fa_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2859 U$$2859/A U$$2871/B VGND VGND VPWR VPWR U$$2859/X sky130_fd_sc_hd__xor2_1
XFILLER_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_801__853 VGND VGND VPWR VPWR _801__853/HI U$$4447/B sky130_fd_sc_hd__conb_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _447_/CLK _426_/D VGND VGND VPWR VPWR _426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_357_ _488_/CLK _357_/D VGND VGND VPWR VPWR _357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_288_ _612_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_80_5 dadda_fa_2_80_5/A dadda_fa_2_80_5/B dadda_fa_2_80_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_2/A dadda_fa_4_80_0/A sky130_fd_sc_hd__fa_1
XFILLER_64_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_73_4 dadda_fa_2_73_4/A dadda_fa_2_73_4/B dadda_fa_2_73_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/CIN dadda_fa_3_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_66_3 dadda_fa_2_66_3/A dadda_fa_2_66_3/B dadda_fa_2_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/B dadda_fa_3_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_69_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_59_2 dadda_fa_2_59_2/A dadda_fa_2_59_2/B dadda_fa_2_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/A dadda_fa_3_59_3/A sky130_fd_sc_hd__fa_2
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 a[12] VGND VGND VPWR VPWR _628_/D sky130_fd_sc_hd__buf_2
Xdadda_fa_5_36_1 dadda_fa_5_36_1/A dadda_fa_5_36_1/B dadda_fa_5_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/B dadda_fa_7_36_0/A sky130_fd_sc_hd__fa_1
XFILLER_37_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_29_0 dadda_fa_5_29_0/A dadda_fa_5_29_0/B dadda_fa_5_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/A dadda_fa_6_29_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_25_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_110_1 dadda_fa_5_110_1/A dadda_fa_5_110_1/B dadda_fa_5_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/B dadda_fa_7_110_0/A sky130_fd_sc_hd__fa_2
XFILLER_118_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$2 _426_/Q _298_/Q VGND VGND VPWR VPWR final_adder.U$$497/B1 final_adder.U$$624/A
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_5_103_0 dadda_fa_5_103_0/A dadda_fa_5_103_0/B dadda_fa_5_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/A dadda_fa_6_103_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput330 _218_/Q VGND VGND VPWR VPWR o[50] sky130_fd_sc_hd__buf_2
XFILLER_134_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput341 _228_/Q VGND VGND VPWR VPWR o[60] sky130_fd_sc_hd__buf_2
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput352 _238_/Q VGND VGND VPWR VPWR o[70] sky130_fd_sc_hd__buf_2
XFILLER_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput363 _248_/Q VGND VGND VPWR VPWR o[80] sky130_fd_sc_hd__buf_2
XFILLER_160_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput374 _258_/Q VGND VGND VPWR VPWR o[90] sky130_fd_sc_hd__buf_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_61_2 U$$2789/X U$$2922/X U$$3055/X VGND VGND VPWR VPWR dadda_fa_2_62_1/A
+ dadda_fa_2_61_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_54_1 U$$1179/X U$$1312/X U$$1445/X VGND VGND VPWR VPWR dadda_fa_2_55_0/CIN
+ dadda_fa_2_54_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_31_0 dadda_fa_4_31_0/A dadda_fa_4_31_0/B dadda_fa_4_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/A dadda_fa_5_31_1/A sky130_fd_sc_hd__fa_1
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_47_0 U$$101/X U$$234/X U$$367/X VGND VGND VPWR VPWR dadda_fa_2_48_1/B
+ dadda_fa_2_47_4/A sky130_fd_sc_hd__fa_2
XFILLER_56_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_211_ _456_/CLK _211_/D VGND VGND VPWR VPWR _211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_83_3 dadda_fa_3_83_3/A dadda_fa_3_83_3/B dadda_fa_3_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/B dadda_fa_4_83_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_2 dadda_fa_3_76_2/A dadda_fa_3_76_2/B dadda_fa_3_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/A dadda_fa_4_76_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_69_1 dadda_fa_3_69_1/A dadda_fa_3_69_1/B dadda_fa_3_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/CIN dadda_fa_4_69_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_46_0 dadda_fa_6_46_0/A dadda_fa_6_46_0/B dadda_fa_6_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_47_0/B dadda_fa_7_46_0/CIN sky130_fd_sc_hd__fa_2
XU$$4003 _563_/Q U$$3977/X _564_/Q U$$3978/X VGND VGND VPWR VPWR U$$4004/A sky130_fd_sc_hd__a22o_1
XU$$4014 U$$4014/A U$$4109/A VGND VGND VPWR VPWR U$$4014/X sky130_fd_sc_hd__xor2_1
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4025 _574_/Q U$$4045/A2 U$$4438/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$4026/A sky130_fd_sc_hd__a22o_1
XU$$4036 U$$4036/A U$$4044/B VGND VGND VPWR VPWR U$$4036/X sky130_fd_sc_hd__xor2_1
XU$$3302 U$$14/A1 U$$3396/A2 _556_/Q U$$3396/B2 VGND VGND VPWR VPWR U$$3303/A sky130_fd_sc_hd__a22o_1
XFILLER_93_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4047 U$$759/A1 U$$4107/A2 U$$759/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4048/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3313 U$$3313/A U$$3413/B VGND VGND VPWR VPWR U$$3313/X sky130_fd_sc_hd__xor2_1
XU$$4058 U$$4058/A U$$4058/B VGND VGND VPWR VPWR U$$4058/X sky130_fd_sc_hd__xor2_1
XU$$4069 _596_/Q U$$4107/A2 U$$98/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4070/A sky130_fd_sc_hd__a22o_1
XU$$3324 U$$4283/A1 U$$3412/A2 U$$4285/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3325/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3335 U$$3335/A U$$3397/B VGND VGND VPWR VPWR U$$3335/X sky130_fd_sc_hd__xor2_1
XU$$3346 _577_/Q U$$3292/X U$$4170/A1 U$$3293/X VGND VGND VPWR VPWR U$$3347/A sky130_fd_sc_hd__a22o_1
XU$$2601 U$$2601/A U$$2603/A VGND VGND VPWR VPWR U$$2601/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2612 U$$2612/A U$$2710/B VGND VGND VPWR VPWR U$$2612/X sky130_fd_sc_hd__xor2_1
XFILLER_34_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_105_2 dadda_fa_4_105_2/A dadda_fa_4_105_2/B dadda_fa_4_105_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/CIN dadda_fa_5_105_1/CIN sky130_fd_sc_hd__fa_1
XU$$3357 U$$3357/A U$$3413/B VGND VGND VPWR VPWR U$$3357/X sky130_fd_sc_hd__xor2_1
XU$$2623 U$$979/A1 U$$2667/A2 U$$979/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2624/A sky130_fd_sc_hd__a22o_1
XFILLER_61_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3368 U$$765/A1 U$$3412/A2 U$$630/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3369/A sky130_fd_sc_hd__a22o_1
XU$$3379 U$$3379/A U$$3403/B VGND VGND VPWR VPWR U$$3379/X sky130_fd_sc_hd__xor2_1
XU$$2634 U$$2634/A U$$2694/B VGND VGND VPWR VPWR U$$2634/X sky130_fd_sc_hd__xor2_1
XFILLER_74_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2645 U$$4289/A1 U$$2667/A2 U$$4289/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2646/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1900 U$$1900/A _643_/Q VGND VGND VPWR VPWR U$$1900/X sky130_fd_sc_hd__xor2_1
XFILLER_46_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1911 U$$952/A1 U$$1785/X U$$952/B1 U$$1786/X VGND VGND VPWR VPWR U$$1912/A sky130_fd_sc_hd__a22o_1
XU$$2656 U$$2656/A U$$2694/B VGND VGND VPWR VPWR U$$2656/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1922 U$$1920/Y _644_/Q U$$1918/A U$$1921/X U$$1918/Y VGND VGND VPWR VPWR U$$1922/X
+ sky130_fd_sc_hd__a32o_4
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2667 U$$3900/A1 U$$2667/A2 U$$3489/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2668/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1933 U$$1933/A U$$1991/B VGND VGND VPWR VPWR U$$1933/X sky130_fd_sc_hd__xor2_1
XU$$2678 U$$2678/A U$$2698/B VGND VGND VPWR VPWR U$$2678/X sky130_fd_sc_hd__xor2_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2689 _591_/Q U$$2607/X U$$4335/A1 U$$2608/X VGND VGND VPWR VPWR U$$2690/A sky130_fd_sc_hd__a22o_1
XFILLER_15_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1944 U$$26/A1 U$$1922/X U$$28/A1 U$$1923/X VGND VGND VPWR VPWR U$$1945/A sky130_fd_sc_hd__a22o_1
XU$$1955 U$$1955/A U$$1991/B VGND VGND VPWR VPWR U$$1955/X sky130_fd_sc_hd__xor2_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1966 U$$48/A1 U$$2048/A2 U$$50/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1967/A sky130_fd_sc_hd__a22o_1
XU$$1977 U$$1977/A U$$1991/B VGND VGND VPWR VPWR U$$1977/X sky130_fd_sc_hd__xor2_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1988 U$$892/A1 U$$2036/A2 U$$892/B1 U$$2036/B2 VGND VGND VPWR VPWR U$$1989/A sky130_fd_sc_hd__a22o_1
XU$$1999 U$$1999/A U$$2021/B VGND VGND VPWR VPWR U$$1999/X sky130_fd_sc_hd__xor2_1
X_409_ _595_/CLK _409_/D VGND VGND VPWR VPWR _409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_119_0 dadda_fa_7_119_0/A dadda_fa_7_119_0/B dadda_fa_7_119_0/CIN VGND
+ VGND VPWR VPWR _544_/D _415_/D sky130_fd_sc_hd__fa_2
XFILLER_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_71_1 dadda_fa_2_71_1/A dadda_fa_2_71_1/B dadda_fa_2_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/CIN dadda_fa_3_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_64_0 dadda_fa_2_64_0/A dadda_fa_2_64_0/B dadda_fa_2_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/B dadda_fa_3_64_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$607 final_adder.U$$734/A final_adder.U$$734/B final_adder.U$$607/B1
+ VGND VGND VPWR VPWR final_adder.U$$735/B sky130_fd_sc_hd__a21o_1
XFILLER_97_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$629 final_adder.U$$7/SUM final_adder.U$$629/B VGND VGND VPWR VPWR
+ hold3/A sky130_fd_sc_hd__xor2_4
XFILLER_111_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$40 U$$40/A1 U$$4/X _569_/Q U$$5/X VGND VGND VPWR VPWR U$$41/A sky130_fd_sc_hd__a22o_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$51 U$$51/A U$$9/B VGND VGND VPWR VPWR U$$51/X sky130_fd_sc_hd__xor2_1
XU$$62 U$$62/A1 U$$4/X U$$64/A1 U$$5/X VGND VGND VPWR VPWR U$$63/A sky130_fd_sc_hd__a22o_1
XU$$73 U$$73/A U$$9/B VGND VGND VPWR VPWR U$$73/X sky130_fd_sc_hd__xor2_1
XU$$84 U$$84/A1 U$$4/X U$$86/A1 U$$5/X VGND VGND VPWR VPWR U$$85/A sky130_fd_sc_hd__a22o_1
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3880 _570_/Q U$$3970/A2 _571_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3881/A sky130_fd_sc_hd__a22o_1
XU$$95 U$$95/A U$$3/A VGND VGND VPWR VPWR U$$95/X sky130_fd_sc_hd__xor2_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3891 U$$3891/A U$$3893/B VGND VGND VPWR VPWR U$$3891/X sky130_fd_sc_hd__xor2_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_93_2 dadda_fa_4_93_2/A dadda_fa_4_93_2/B dadda_fa_4_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/CIN dadda_fa_5_93_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_86_1 dadda_fa_4_86_1/A dadda_fa_4_86_1/B dadda_fa_4_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/B dadda_fa_5_86_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_63_0 dadda_fa_7_63_0/A dadda_fa_7_63_0/B dadda_fa_7_63_0/CIN VGND VGND
+ VPWR VPWR _488_/D _359_/D sky130_fd_sc_hd__fa_1
XFILLER_133_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_79_0 dadda_fa_4_79_0/A dadda_fa_4_79_0/B dadda_fa_4_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/A dadda_fa_5_79_1/A sky130_fd_sc_hd__fa_2
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1207 U$$1207/A U$$1232/A VGND VGND VPWR VPWR U$$1207/X sky130_fd_sc_hd__xor2_1
XU$$1218 _609_/Q U$$1218/A2 _610_/Q U$$1218/B2 VGND VGND VPWR VPWR U$$1219/A sky130_fd_sc_hd__a22o_1
XFILLER_16_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1229 U$$1229/A _633_/Q VGND VGND VPWR VPWR U$$1229/X sky130_fd_sc_hd__xor2_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_81_0 dadda_fa_3_81_0/A dadda_fa_3_81_0/B dadda_fa_3_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/B dadda_fa_4_81_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_113_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3110 U$$96/A1 U$$3018/X _597_/Q U$$3019/X VGND VGND VPWR VPWR U$$3111/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_0 input141/X dadda_fa_4_110_0/B dadda_fa_4_110_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_111_0/A dadda_fa_5_110_1/A sky130_fd_sc_hd__fa_1
XU$$3121 U$$3121/A _661_/Q VGND VGND VPWR VPWR U$$3121/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_43_5 dadda_fa_2_43_5/A dadda_fa_2_43_5/B dadda_fa_2_43_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_2/A dadda_fa_4_43_0/A sky130_fd_sc_hd__fa_2
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3132 U$$4502/A1 U$$3018/X U$$4504/A1 U$$3019/X VGND VGND VPWR VPWR U$$3133/A sky130_fd_sc_hd__a22o_1
XU$$3143 U$$3143/A _661_/Q VGND VGND VPWR VPWR U$$3143/X sky130_fd_sc_hd__xor2_1
XU$$3154 U$$3270/B U$$3154/B VGND VGND VPWR VPWR U$$3154/X sky130_fd_sc_hd__and2_1
Xdadda_fa_2_36_4 U$$2340/X U$$2473/X U$$2533/B VGND VGND VPWR VPWR dadda_fa_3_37_1/CIN
+ dadda_fa_3_36_3/CIN sky130_fd_sc_hd__fa_1
XU$$3165 U$$14/A1 U$$3243/A2 _556_/Q U$$3243/B2 VGND VGND VPWR VPWR U$$3166/A sky130_fd_sc_hd__a22o_1
XFILLER_62_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2420 U$$2420/A U$$2432/B VGND VGND VPWR VPWR U$$2420/X sky130_fd_sc_hd__xor2_1
XFILLER_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2431 U$$924/A1 U$$2463/A2 U$$926/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2432/A sky130_fd_sc_hd__a22o_1
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3176 U$$3176/A U$$3224/B VGND VGND VPWR VPWR U$$3176/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2442 U$$2442/A U$$2464/B VGND VGND VPWR VPWR U$$2442/X sky130_fd_sc_hd__xor2_1
XU$$3187 U$$4283/A1 U$$3241/A2 U$$4285/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3188/A
+ sky130_fd_sc_hd__a22o_1
XU$$2453 _610_/Q U$$2463/A2 U$$4510/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2454/A sky130_fd_sc_hd__a22o_1
XU$$3198 U$$3198/A U$$3224/B VGND VGND VPWR VPWR U$$3198/X sky130_fd_sc_hd__xor2_1
XU$$2464 U$$2464/A U$$2464/B VGND VGND VPWR VPWR U$$2464/X sky130_fd_sc_hd__xor2_1
XFILLER_50_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1730 U$$771/A1 U$$1734/A2 U$$771/B1 U$$1734/B2 VGND VGND VPWR VPWR U$$1731/A sky130_fd_sc_hd__a22o_1
XU$$2475 U$$2475/A U$$2533/B VGND VGND VPWR VPWR U$$2475/X sky130_fd_sc_hd__xor2_1
XFILLER_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1741 U$$1741/A U$$1781/A VGND VGND VPWR VPWR U$$1741/X sky130_fd_sc_hd__xor2_1
XFILLER_62_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2486 U$$979/A1 U$$2534/A2 U$$979/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2487/A sky130_fd_sc_hd__a22o_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1752 U$$928/B1 U$$1648/X _603_/Q U$$1649/X VGND VGND VPWR VPWR U$$1753/A sky130_fd_sc_hd__a22o_1
XU$$2497 U$$2497/A U$$2533/B VGND VGND VPWR VPWR U$$2497/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1763 U$$1763/A U$$1781/A VGND VGND VPWR VPWR U$$1763/X sky130_fd_sc_hd__xor2_1
XFILLER_188_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1774 U$$4514/A1 U$$1648/X U$$952/B1 U$$1649/X VGND VGND VPWR VPWR U$$1775/A sky130_fd_sc_hd__a22o_1
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1785 U$$1783/Y _642_/Q U$$1781/A U$$1784/X U$$1781/Y VGND VGND VPWR VPWR U$$1785/X
+ sky130_fd_sc_hd__a32o_4
XU$$1796 U$$1796/A U$$1918/A VGND VGND VPWR VPWR U$$1796/X sky130_fd_sc_hd__xor2_1
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_96_0 dadda_fa_5_96_0/A dadda_fa_5_96_0/B dadda_fa_5_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/A dadda_fa_6_96_0/CIN sky130_fd_sc_hd__fa_1
Xinput40 a[45] VGND VGND VPWR VPWR _661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 a[55] VGND VGND VPWR VPWR _671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput62 a[7] VGND VGND VPWR VPWR _623_/D sky130_fd_sc_hd__clkbuf_4
Xinput73 b[17] VGND VGND VPWR VPWR _569_/D sky130_fd_sc_hd__clkbuf_4
Xinput84 b[27] VGND VGND VPWR VPWR _579_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput95 b[37] VGND VGND VPWR VPWR _589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$415 final_adder.U$$332/B final_adder.U$$670/B final_adder.U$$281/X
+ VGND VGND VPWR VPWR final_adder.U$$674/B sky130_fd_sc_hd__a21o_1
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater630 _606_/Q VGND VGND VPWR VPWR U$$938/A1 sky130_fd_sc_hd__buf_12
XFILLER_57_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$437 final_adder.U$$260/B final_adder.U$$630/B final_adder.U$$137/X
+ VGND VGND VPWR VPWR final_adder.U$$632/B sky130_fd_sc_hd__a21o_1
Xrepeater641 _601_/Q VGND VGND VPWR VPWR U$$654/A1 sky130_fd_sc_hd__buf_12
XFILLER_123_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater652 U$$96/A1 VGND VGND VPWR VPWR U$$94/B1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$459 final_adder.U$$282/B final_adder.U$$674/B final_adder.U$$181/X
+ VGND VGND VPWR VPWR final_adder.U$$676/B sky130_fd_sc_hd__a21o_1
Xrepeater663 _592_/Q VGND VGND VPWR VPWR U$$4335/A1 sky130_fd_sc_hd__buf_12
Xrepeater674 _588_/Q VGND VGND VPWR VPWR U$$765/A1 sky130_fd_sc_hd__buf_12
XU$$309 U$$309/A U$$391/B VGND VGND VPWR VPWR U$$309/X sky130_fd_sc_hd__xor2_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater685 _584_/Q VGND VGND VPWR VPWR U$$72/A1 sky130_fd_sc_hd__buf_12
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater696 U$$4446/A1 VGND VGND VPWR VPWR U$$62/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_105_1 U$$4074/X U$$4207/X U$$4340/X VGND VGND VPWR VPWR dadda_fa_4_106_0/CIN
+ dadda_fa_4_105_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_126_0 U$$4515/X input158/X dadda_fa_6_126_0/CIN VGND VGND VPWR VPWR dadda_fa_7_127_0/B
+ dadda_fa_7_126_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_69_4 U$$2007/X U$$2140/X U$$2273/X VGND VGND VPWR VPWR dadda_fa_1_70_7/B
+ dadda_fa_2_69_0/A sky130_fd_sc_hd__fa_2
XFILLER_75_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_46_3 dadda_fa_3_46_3/A dadda_fa_3_46_3/B dadda_fa_3_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/B dadda_fa_4_46_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$810 U$$810/A _627_/Q VGND VGND VPWR VPWR U$$810/X sky130_fd_sc_hd__xor2_1
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_674_ _679_/CLK _674_/D VGND VGND VPWR VPWR _674_/Q sky130_fd_sc_hd__dfxtp_2
XU$$821 _627_/Q VGND VGND VPWR VPWR U$$821/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_3_39_2 dadda_fa_3_39_2/A dadda_fa_3_39_2/B dadda_fa_3_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/A dadda_fa_4_39_2/B sky130_fd_sc_hd__fa_2
XU$$832 U$$8/B1 U$$928/A2 U$$971/A1 U$$928/B2 VGND VGND VPWR VPWR U$$833/A sky130_fd_sc_hd__a22o_1
XU$$843 U$$843/A U$$959/A VGND VGND VPWR VPWR U$$843/X sky130_fd_sc_hd__xor2_1
XFILLER_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$854 U$$32/A1 U$$910/A2 U$$34/A1 U$$910/B2 VGND VGND VPWR VPWR U$$855/A sky130_fd_sc_hd__a22o_1
XU$$865 U$$865/A U$$959/A VGND VGND VPWR VPWR U$$865/X sky130_fd_sc_hd__xor2_1
XU$$1004 U$$1004/A U$$980/B VGND VGND VPWR VPWR U$$1004/X sky130_fd_sc_hd__xor2_1
XU$$1015 U$$878/A1 U$$999/A2 U$$58/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1016/A sky130_fd_sc_hd__a22o_1
XU$$876 U$$876/A1 U$$910/A2 U$$878/A1 U$$910/B2 VGND VGND VPWR VPWR U$$877/A sky130_fd_sc_hd__a22o_1
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1026 U$$1026/A U$$980/B VGND VGND VPWR VPWR U$$1026/X sky130_fd_sc_hd__xor2_1
XU$$887 U$$887/A U$$959/A VGND VGND VPWR VPWR U$$887/X sky130_fd_sc_hd__xor2_1
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1037 U$$78/A1 U$$1093/A2 U$$80/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1038/A sky130_fd_sc_hd__a22o_1
XU$$898 U$$76/A1 U$$910/A2 U$$76/B1 U$$910/B2 VGND VGND VPWR VPWR U$$899/A sky130_fd_sc_hd__a22o_1
XU$$1048 U$$1048/A U$$980/B VGND VGND VPWR VPWR U$$1048/X sky130_fd_sc_hd__xor2_1
XU$$1059 U$$785/A1 U$$1093/A2 U$$924/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1060/A sky130_fd_sc_hd__a22o_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_41_2 U$$2350/X U$$2483/X U$$2616/X VGND VGND VPWR VPWR dadda_fa_3_42_1/A
+ dadda_fa_3_41_3/A sky130_fd_sc_hd__fa_1
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_34_1 U$$740/X U$$873/X U$$1006/X VGND VGND VPWR VPWR dadda_fa_3_35_0/CIN
+ dadda_fa_3_34_2/CIN sky130_fd_sc_hd__fa_1
XU$$2250 U$$4442/A1 U$$2270/A2 U$$4170/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2251/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_0 U$$694/X input151/X dadda_fa_5_11_0/CIN VGND VGND VPWR VPWR dadda_fa_6_12_0/A
+ dadda_fa_6_11_0/CIN sky130_fd_sc_hd__fa_1
XU$$2261 U$$2261/A U$$2327/B VGND VGND VPWR VPWR U$$2261/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_27_0 U$$61/X U$$194/X U$$327/X VGND VGND VPWR VPWR dadda_fa_3_28_2/A dadda_fa_3_27_3/B
+ sky130_fd_sc_hd__fa_2
XU$$2272 U$$80/A1 U$$2316/A2 U$$630/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2273/A sky130_fd_sc_hd__a22o_1
XFILLER_90_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2283 U$$2283/A U$$2327/B VGND VGND VPWR VPWR U$$2283/X sky130_fd_sc_hd__xor2_1
XU$$2294 U$$4486/A1 U$$2316/A2 U$$787/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2295/A
+ sky130_fd_sc_hd__a22o_1
XU$$1560 U$$1560/A U$$1580/B VGND VGND VPWR VPWR U$$1560/X sky130_fd_sc_hd__xor2_1
XU$$1571 U$$3900/A1 U$$1605/A2 U$$3489/B1 U$$1605/B2 VGND VGND VPWR VPWR U$$1572/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1582 U$$1582/A U$$1643/A VGND VGND VPWR VPWR U$$1582/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1593 U$$86/A1 U$$1605/A2 U$$88/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1594/A sky130_fd_sc_hd__a22o_1
XFILLER_33_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_86_4 U$$3105/X U$$3238/X U$$3371/X VGND VGND VPWR VPWR dadda_fa_2_87_4/A
+ dadda_fa_2_86_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_79_3 U$$2293/X U$$2426/X U$$2559/X VGND VGND VPWR VPWR dadda_fa_2_80_1/B
+ dadda_fa_2_79_4/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_56_2 dadda_fa_4_56_2/A dadda_fa_4_56_2/B dadda_fa_4_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/CIN dadda_fa_5_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$201 final_adder.U$$695/A final_adder.U$$567/B1 final_adder.U$$201/B1
+ VGND VGND VPWR VPWR final_adder.U$$201/X sky130_fd_sc_hd__a21o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$212 final_adder.U$$707/A final_adder.U$$706/A VGND VGND VPWR VPWR
+ final_adder.U$$298/B sky130_fd_sc_hd__and2_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$223 final_adder.U$$717/A final_adder.U$$589/B1 final_adder.U$$223/B1
+ VGND VGND VPWR VPWR final_adder.U$$223/X sky130_fd_sc_hd__a21o_1
XFILLER_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_49_1 dadda_fa_4_49_1/A dadda_fa_4_49_1/B dadda_fa_4_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/B dadda_fa_5_49_1/B sky130_fd_sc_hd__fa_1
XFILLER_100_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$234 final_adder.U$$729/A final_adder.U$$728/A VGND VGND VPWR VPWR
+ final_adder.U$$308/A sky130_fd_sc_hd__and2_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$245 final_adder.U$$739/A final_adder.U$$611/B1 final_adder.U$$245/B1
+ VGND VGND VPWR VPWR final_adder.U$$245/X sky130_fd_sc_hd__a21o_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_26_0 dadda_fa_7_26_0/A dadda_fa_7_26_0/B dadda_fa_7_26_0/CIN VGND VGND
+ VPWR VPWR _451_/D _322_/D sky130_fd_sc_hd__fa_2
Xrepeater460 U$$4252/X VGND VGND VPWR VPWR U$$4381/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$267 final_adder.U$$266/A final_adder.U$$149/X final_adder.U$$151/X
+ VGND VGND VPWR VPWR final_adder.U$$267/X sky130_fd_sc_hd__a21o_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$106 U$$928/A1 U$$4/X U$$930/A1 U$$5/X VGND VGND VPWR VPWR U$$107/A sky130_fd_sc_hd__a22o_1
Xrepeater471 U$$3567/X VGND VGND VPWR VPWR U$$3668/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$278 final_adder.U$$278/A final_adder.U$$278/B VGND VGND VPWR VPWR
+ final_adder.U$$330/A sky130_fd_sc_hd__and2_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$117 U$$117/A U$$89/B VGND VGND VPWR VPWR U$$117/X sky130_fd_sc_hd__xor2_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater482 U$$2826/B2 VGND VGND VPWR VPWR U$$2834/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$289 final_adder.U$$288/A final_adder.U$$193/X final_adder.U$$195/X
+ VGND VGND VPWR VPWR final_adder.U$$289/X sky130_fd_sc_hd__a21o_1
Xrepeater493 U$$2197/X VGND VGND VPWR VPWR U$$2316/B2 sky130_fd_sc_hd__buf_12
XU$$128 U$$950/A1 U$$4/X U$$952/A1 U$$5/X VGND VGND VPWR VPWR U$$129/A sky130_fd_sc_hd__a22o_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$139 U$$274/A VGND VGND VPWR VPWR U$$139/Y sky130_fd_sc_hd__inv_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_390_ _535_/CLK _390_/D VGND VGND VPWR VPWR _390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput230 c[76] VGND VGND VPWR VPWR input230/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_3_51_1 dadda_fa_3_51_1/A dadda_fa_3_51_1/B dadda_fa_3_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/CIN dadda_fa_4_51_2/A sky130_fd_sc_hd__fa_1
Xinput241 c[86] VGND VGND VPWR VPWR input241/X sky130_fd_sc_hd__buf_2
Xinput252 c[96] VGND VGND VPWR VPWR input252/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_67_1 U$$540/X U$$673/X U$$806/X VGND VGND VPWR VPWR dadda_fa_1_68_5/CIN
+ dadda_fa_1_67_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_44_0 dadda_fa_3_44_0/A dadda_fa_3_44_0/B dadda_fa_3_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/B dadda_fa_4_44_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$640 U$$92/A1 U$$682/A2 U$$92/B1 U$$553/X VGND VGND VPWR VPWR U$$641/A sky130_fd_sc_hd__a22o_1
X_657_ _667_/CLK _657_/D VGND VGND VPWR VPWR _657_/Q sky130_fd_sc_hd__dfxtp_4
XU$$651 U$$651/A _625_/Q VGND VGND VPWR VPWR U$$651/X sky130_fd_sc_hd__xor2_1
XU$$662 U$$799/A1 U$$682/A2 U$$938/A1 U$$553/X VGND VGND VPWR VPWR U$$663/A sky130_fd_sc_hd__a22o_1
XU$$673 U$$673/A _625_/Q VGND VGND VPWR VPWR U$$673/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$684 _625_/Q VGND VGND VPWR VPWR U$$684/Y sky130_fd_sc_hd__inv_1
XFILLER_189_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$695 U$$8/B1 U$$785/A2 U$$12/A1 U$$785/B2 VGND VGND VPWR VPWR U$$696/A sky130_fd_sc_hd__a22o_1
X_588_ _601_/CLK _588_/D VGND VGND VPWR VPWR _588_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_101_0 dadda_fa_7_101_0/A dadda_fa_7_101_0/B dadda_fa_7_101_0/CIN VGND
+ VGND VPWR VPWR _526_/D _397_/D sky130_fd_sc_hd__fa_2
XFILLER_157_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_96_3 U$$3657/X U$$3790/X U$$3923/X VGND VGND VPWR VPWR dadda_fa_3_97_1/B
+ dadda_fa_3_96_3/B sky130_fd_sc_hd__fa_2
XFILLER_67_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_89_2 U$$4175/X U$$4308/X U$$4441/X VGND VGND VPWR VPWR dadda_fa_3_90_1/A
+ dadda_fa_3_89_3/A sky130_fd_sc_hd__fa_2
XFILLER_126_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_66_1 dadda_fa_5_66_1/A dadda_fa_5_66_1/B dadda_fa_5_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/B dadda_fa_7_66_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_59_0 dadda_fa_5_59_0/A dadda_fa_5_59_0/B dadda_fa_5_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/A dadda_fa_6_59_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_58_8 dadda_fa_1_58_8/A dadda_fa_1_58_8/B dadda_fa_1_58_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_3/A dadda_fa_3_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_105_0 U$$2876/Y U$$3010/X U$$3143/X VGND VGND VPWR VPWR dadda_fa_3_106_3/A
+ dadda_fa_3_105_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2080 U$$2080/A U$$2186/B VGND VGND VPWR VPWR U$$2080/X sky130_fd_sc_hd__xor2_1
XU$$2091 U$$4283/A1 U$$2117/A2 U$$4285/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1390 U$$20/A1 U$$1474/A2 _559_/Q U$$1466/B2 VGND VGND VPWR VPWR U$$1391/A sky130_fd_sc_hd__a22o_1
XFILLER_182_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_91_2 U$$2716/X U$$2849/X U$$2982/X VGND VGND VPWR VPWR dadda_fa_2_92_5/A
+ dadda_fa_3_91_0/A sky130_fd_sc_hd__fa_2
XFILLER_163_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_84_1 U$$1771/X U$$1904/X U$$2037/X VGND VGND VPWR VPWR dadda_fa_2_85_2/B
+ dadda_fa_2_84_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_712__764 VGND VGND VPWR VPWR _712__764/HI U$$1102/A1 sky130_fd_sc_hd__conb_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_61_0 dadda_fa_4_61_0/A dadda_fa_4_61_0/B dadda_fa_4_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/A dadda_fa_5_61_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_0 U$$1358/X U$$1491/X U$$1624/X VGND VGND VPWR VPWR dadda_fa_2_78_0/B
+ dadda_fa_2_77_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_104_2 U$$3540/X U$$3673/X VGND VGND VPWR VPWR dadda_fa_3_105_3/B dadda_fa_4_104_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3709 U$$969/A1 U$$3783/A2 U$$12/A1 U$$3783/B2 VGND VGND VPWR VPWR U$$3710/A sky130_fd_sc_hd__a22o_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ _518_/CLK _511_/D VGND VGND VPWR VPWR _511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _455_/CLK _442_/D VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_373_ _500_/CLK _373_/D VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_99_1 dadda_fa_3_99_1/A dadda_fa_3_99_1/B dadda_fa_3_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_0/CIN dadda_fa_4_99_2/A sky130_fd_sc_hd__fa_2
XFILLER_86_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_76_0 dadda_fa_6_76_0/A dadda_fa_6_76_0/B dadda_fa_6_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_77_0/B dadda_fa_7_76_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_181_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_702__922 VGND VGND VPWR VPWR _702__922/HI _702__922/LO sky130_fd_sc_hd__conb_1
XU$$470 U$$470/A _623_/Q VGND VGND VPWR VPWR U$$470/X sky130_fd_sc_hd__xor2_1
XFILLER_45_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$481 U$$70/A1 U$$545/A2 U$$70/B1 U$$416/X VGND VGND VPWR VPWR U$$482/A sky130_fd_sc_hd__a22o_1
XU$$492 U$$492/A U$$547/A VGND VGND VPWR VPWR U$$492/X sky130_fd_sc_hd__xor2_1
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_94_0 U$$2722/X U$$2855/X U$$2988/X VGND VGND VPWR VPWR dadda_fa_3_95_0/B
+ dadda_fa_3_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_7 dadda_fa_1_70_7/A dadda_fa_1_70_7/B dadda_fa_1_70_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/CIN dadda_fa_2_70_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_6 dadda_fa_1_63_6/A dadda_fa_1_63_6/B dadda_fa_1_63_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/B dadda_fa_2_63_5/B sky130_fd_sc_hd__fa_1
XFILLER_189_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_56_5 U$$3178/X U$$3311/X U$$3444/X VGND VGND VPWR VPWR dadda_fa_2_57_2/A
+ dadda_fa_2_56_5/A sky130_fd_sc_hd__fa_1
XFILLER_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_49_4 U$$1701/X U$$1834/X U$$1967/X VGND VGND VPWR VPWR dadda_fa_2_50_2/A
+ dadda_fa_2_49_5/A sky130_fd_sc_hd__fa_1
XFILLER_55_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_2 dadda_fa_4_19_2/A dadda_fa_4_19_2/B dadda_ha_3_19_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/CIN dadda_fa_5_19_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_93_0 dadda_fa_7_93_0/A dadda_fa_7_93_0/B dadda_fa_7_93_0/CIN VGND VGND
+ VPWR VPWR _518_/D _389_/D sky130_fd_sc_hd__fa_1
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4207 U$$4207/A _677_/Q VGND VGND VPWR VPWR U$$4207/X sky130_fd_sc_hd__xor2_1
XU$$4218 U$$4492/A1 U$$4114/X U$$4494/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4219/A
+ sky130_fd_sc_hd__a22o_1
XU$$4229 U$$4229/A U$$4246/A VGND VGND VPWR VPWR U$$4229/X sky130_fd_sc_hd__xor2_1
XFILLER_120_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3506 U$$3506/A _667_/Q VGND VGND VPWR VPWR U$$3506/X sky130_fd_sc_hd__xor2_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3517 U$$4476/A1 U$$3545/A2 U$$94/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3518/A sky130_fd_sc_hd__a22o_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3528 U$$3528/A _667_/Q VGND VGND VPWR VPWR U$$3528/X sky130_fd_sc_hd__xor2_1
XFILLER_105_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3539 _605_/Q U$$3429/X U$$4500/A1 U$$3430/X VGND VGND VPWR VPWR U$$3540/A sky130_fd_sc_hd__a22o_1
XFILLER_74_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2805 U$$2805/A U$$2839/B VGND VGND VPWR VPWR U$$2805/X sky130_fd_sc_hd__xor2_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2816 U$$2953/A1 U$$2868/A2 U$$76/B1 U$$2834/B2 VGND VGND VPWR VPWR U$$2817/A sky130_fd_sc_hd__a22o_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2827 U$$2827/A U$$2839/B VGND VGND VPWR VPWR U$$2827/X sky130_fd_sc_hd__xor2_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2838 _597_/Q U$$2868/A2 U$$4484/A1 U$$2745/X VGND VGND VPWR VPWR U$$2839/A sky130_fd_sc_hd__a22o_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2849 U$$2849/A U$$2871/B VGND VGND VPWR VPWR U$$2849/X sky130_fd_sc_hd__xor2_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_2 U$$847/X U$$980/X U$$1113/X VGND VGND VPWR VPWR dadda_fa_4_22_1/A
+ dadda_fa_4_21_2/B sky130_fd_sc_hd__fa_2
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_840__892 VGND VGND VPWR VPWR _840__892/HI U$$6/A1 sky130_fd_sc_hd__conb_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_425_ _425_/CLK _425_/D VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_356_ _488_/CLK _356_/D VGND VGND VPWR VPWR _356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_287_ _612_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_73_5 dadda_fa_2_73_5/A dadda_fa_2_73_5/B dadda_fa_2_73_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_2/A dadda_fa_4_73_0/A sky130_fd_sc_hd__fa_2
XFILLER_151_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_66_4 dadda_fa_2_66_4/A dadda_fa_2_66_4/B dadda_fa_2_66_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/CIN dadda_fa_3_66_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_59_3 dadda_fa_2_59_3/A dadda_fa_2_59_3/B dadda_fa_2_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/B dadda_fa_3_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 a[13] VGND VGND VPWR VPWR _629_/D sky130_fd_sc_hd__buf_2
XFILLER_7_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_29_1 dadda_fa_5_29_1/A dadda_fa_5_29_1/B dadda_fa_5_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/B dadda_fa_7_29_0/A sky130_fd_sc_hd__fa_2
XFILLER_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$3 _427_/Q _299_/Q VGND VGND VPWR VPWR final_adder.U$$3/COUT final_adder.U$$625/A
+ sky130_fd_sc_hd__ha_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_103_1 dadda_fa_5_103_1/A dadda_fa_5_103_1/B dadda_fa_5_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/B dadda_fa_7_103_0/A sky130_fd_sc_hd__fa_2
XFILLER_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput320 _209_/Q VGND VGND VPWR VPWR o[41] sky130_fd_sc_hd__buf_2
XFILLER_156_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput331 _219_/Q VGND VGND VPWR VPWR o[51] sky130_fd_sc_hd__buf_2
Xoutput342 _229_/Q VGND VGND VPWR VPWR o[61] sky130_fd_sc_hd__buf_2
Xoutput353 _239_/Q VGND VGND VPWR VPWR o[71] sky130_fd_sc_hd__buf_2
Xoutput364 _249_/Q VGND VGND VPWR VPWR o[81] sky130_fd_sc_hd__buf_2
XFILLER_126_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput375 _259_/Q VGND VGND VPWR VPWR o[91] sky130_fd_sc_hd__buf_2
XFILLER_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_783__835 VGND VGND VPWR VPWR _783__835/HI U$$4411/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_61_3 U$$3188/X U$$3321/X U$$3454/X VGND VGND VPWR VPWR dadda_fa_2_62_1/B
+ dadda_fa_2_61_4/B sky130_fd_sc_hd__fa_1
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_2 U$$1578/X U$$1711/X U$$1844/X VGND VGND VPWR VPWR dadda_fa_2_55_1/A
+ dadda_fa_2_54_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_31_1 dadda_fa_4_31_1/A dadda_fa_4_31_1/B dadda_fa_4_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/B dadda_fa_5_31_1/B sky130_fd_sc_hd__fa_2
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_1 U$$500/X U$$633/X U$$766/X VGND VGND VPWR VPWR dadda_fa_2_48_1/CIN
+ dadda_fa_2_47_4/B sky130_fd_sc_hd__fa_2
X_824__876 VGND VGND VPWR VPWR _824__876/HI U$$4493/B sky130_fd_sc_hd__conb_1
Xdadda_fa_4_24_0 dadda_fa_4_24_0/A dadda_fa_4_24_0/B dadda_fa_4_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/A dadda_fa_5_24_1/A sky130_fd_sc_hd__fa_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_210_ _329_/CLK _210_/D VGND VGND VPWR VPWR _210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_718__770 VGND VGND VPWR VPWR _718__770/HI U$$143/A1 sky130_fd_sc_hd__conb_1
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_76_3 dadda_fa_3_76_3/A dadda_fa_3_76_3/B dadda_fa_3_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/B dadda_fa_4_76_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_69_2 dadda_fa_3_69_2/A dadda_fa_3_69_2/B dadda_fa_3_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/A dadda_fa_4_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_104_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4004 U$$4004/A U$$4058/B VGND VGND VPWR VPWR U$$4004/X sky130_fd_sc_hd__xor2_1
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4015 _569_/Q U$$4107/A2 _570_/Q U$$4107/B2 VGND VGND VPWR VPWR U$$4016/A sky130_fd_sc_hd__a22o_1
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4026 U$$4026/A U$$4044/B VGND VGND VPWR VPWR U$$4026/X sky130_fd_sc_hd__xor2_1
XU$$4037 _580_/Q U$$3977/X _581_/Q U$$3978/X VGND VGND VPWR VPWR U$$4038/A sky130_fd_sc_hd__a22o_1
XFILLER_120_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_39_0 dadda_fa_6_39_0/A dadda_fa_6_39_0/B dadda_fa_6_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_40_0/B dadda_fa_7_39_0/CIN sky130_fd_sc_hd__fa_1
XU$$3303 U$$3303/A U$$3397/B VGND VGND VPWR VPWR U$$3303/X sky130_fd_sc_hd__xor2_1
XU$$4048 U$$4048/A U$$4109/A VGND VGND VPWR VPWR U$$4048/X sky130_fd_sc_hd__xor2_1
XFILLER_59_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3314 U$$4273/A1 U$$3396/A2 _562_/Q U$$3396/B2 VGND VGND VPWR VPWR U$$3315/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4059 U$$771/A1 U$$4107/A2 U$$4335/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4060/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3325 U$$3325/A U$$3397/B VGND VGND VPWR VPWR U$$3325/X sky130_fd_sc_hd__xor2_1
XU$$3336 U$$4156/B1 U$$3396/A2 _573_/Q U$$3396/B2 VGND VGND VPWR VPWR U$$3337/A sky130_fd_sc_hd__a22o_1
XU$$3347 U$$3347/A U$$3403/B VGND VGND VPWR VPWR U$$3347/X sky130_fd_sc_hd__xor2_1
XU$$2602 U$$2603/A VGND VGND VPWR VPWR U$$2602/Y sky130_fd_sc_hd__inv_1
XFILLER_46_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2613 U$$8/B1 U$$2729/A2 U$$12/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2614/A sky130_fd_sc_hd__a22o_1
XU$$3358 U$$892/A1 U$$3396/A2 U$$892/B1 U$$3396/B2 VGND VGND VPWR VPWR U$$3359/A sky130_fd_sc_hd__a22o_1
XU$$2624 U$$2624/A U$$2694/B VGND VGND VPWR VPWR U$$2624/X sky130_fd_sc_hd__xor2_1
XU$$3369 U$$3369/A U$$3413/B VGND VGND VPWR VPWR U$$3369/X sky130_fd_sc_hd__xor2_1
XU$$2635 _564_/Q U$$2667/A2 _565_/Q U$$2667/B2 VGND VGND VPWR VPWR U$$2636/A sky130_fd_sc_hd__a22o_1
XFILLER_34_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1901 _608_/Q U$$1903/A2 _609_/Q U$$1903/B2 VGND VGND VPWR VPWR U$$1902/A sky130_fd_sc_hd__a22o_1
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2646 U$$2646/A U$$2694/B VGND VGND VPWR VPWR U$$2646/X sky130_fd_sc_hd__xor2_1
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1912 U$$1912/A _643_/Q VGND VGND VPWR VPWR U$$1912/X sky130_fd_sc_hd__xor2_1
XU$$2657 U$$876/A1 U$$2667/A2 U$$878/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2658/A sky130_fd_sc_hd__a22o_1
XU$$1923 U$$1921/B U$$1918/A _644_/Q U$$1918/Y VGND VGND VPWR VPWR U$$1923/X sky130_fd_sc_hd__a22o_4
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2668 U$$2668/A U$$2694/B VGND VGND VPWR VPWR U$$2668/X sky130_fd_sc_hd__xor2_1
XU$$2679 _586_/Q U$$2607/X _587_/Q U$$2608/X VGND VGND VPWR VPWR U$$2680/A sky130_fd_sc_hd__a22o_1
XFILLER_178_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1934 U$$14/B1 U$$2048/A2 U$$4265/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$1935/A sky130_fd_sc_hd__a22o_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1945 U$$1945/A U$$2021/B VGND VGND VPWR VPWR U$$1945/X sky130_fd_sc_hd__xor2_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1956 U$$4285/A1 U$$2036/A2 U$$3191/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1957/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1967 U$$1967/A U$$1991/B VGND VGND VPWR VPWR U$$1967/X sky130_fd_sc_hd__xor2_1
XU$$1978 U$$4170/A1 U$$2036/A2 U$$3624/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1979/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _594_/CLK _408_/D VGND VGND VPWR VPWR _408_/Q sky130_fd_sc_hd__dfxtp_2
XU$$1989 U$$1989/A U$$2023/B VGND VGND VPWR VPWR U$$1989/X sky130_fd_sc_hd__xor2_1
XFILLER_186_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_339_ _339_/CLK _339_/D VGND VGND VPWR VPWR _339_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_767__819 VGND VGND VPWR VPWR _767__819/HI U$$4385/A sky130_fd_sc_hd__conb_1
XFILLER_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_71_2 dadda_fa_2_71_2/A dadda_fa_2_71_2/B dadda_fa_2_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/A dadda_fa_3_71_3/A sky130_fd_sc_hd__fa_2
XFILLER_155_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_64_1 dadda_fa_2_64_1/A dadda_fa_2_64_1/B dadda_fa_2_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/CIN dadda_fa_3_64_2/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$619 final_adder.U$$746/A final_adder.U$$746/B final_adder.U$$619/B1
+ VGND VGND VPWR VPWR final_adder.U$$747/B sky130_fd_sc_hd__a21o_1
XFILLER_38_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_41_0 dadda_fa_5_41_0/A dadda_fa_5_41_0/B dadda_fa_5_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/A dadda_fa_6_41_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_57_0 dadda_fa_2_57_0/A dadda_fa_2_57_0/B dadda_fa_2_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/B dadda_fa_3_57_2/B sky130_fd_sc_hd__fa_2
XFILLER_116_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$30 U$$30/A1 U$$4/X U$$30/B1 U$$5/X VGND VGND VPWR VPWR U$$31/A sky130_fd_sc_hd__a22o_1
XU$$41 U$$41/A U$$3/A VGND VGND VPWR VPWR U$$41/X sky130_fd_sc_hd__xor2_1
XU$$52 U$$52/A1 U$$4/X U$$54/A1 U$$5/X VGND VGND VPWR VPWR U$$53/A sky130_fd_sc_hd__a22o_1
XU$$63 U$$63/A U$$89/B VGND VGND VPWR VPWR U$$63/X sky130_fd_sc_hd__xor2_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$74 U$$74/A1 U$$4/X U$$76/A1 U$$5/X VGND VGND VPWR VPWR U$$75/A sky130_fd_sc_hd__a22o_1
XU$$3870 _565_/Q U$$3840/X U$$4283/A1 U$$3841/X VGND VGND VPWR VPWR U$$3871/A sky130_fd_sc_hd__a22o_1
XU$$85 U$$85/A U$$9/B VGND VGND VPWR VPWR U$$85/X sky130_fd_sc_hd__xor2_2
XU$$3881 U$$3881/A U$$3969/B VGND VGND VPWR VPWR U$$3881/X sky130_fd_sc_hd__xor2_1
XU$$96 U$$96/A1 U$$4/X U$$96/B1 U$$5/X VGND VGND VPWR VPWR U$$97/A sky130_fd_sc_hd__a22o_1
XFILLER_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3892 U$$56/A1 U$$3912/A2 U$$4442/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3893/A sky130_fd_sc_hd__a22o_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_86_2 dadda_fa_4_86_2/A dadda_fa_4_86_2/B dadda_fa_4_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/CIN dadda_fa_5_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_79_1 dadda_fa_4_79_1/A dadda_fa_4_79_1/B dadda_fa_4_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/B dadda_fa_5_79_1/B sky130_fd_sc_hd__fa_1
XFILLER_115_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_56_0 dadda_fa_7_56_0/A dadda_fa_7_56_0/B dadda_fa_7_56_0/CIN VGND VGND
+ VPWR VPWR _481_/D _352_/D sky130_fd_sc_hd__fa_1
XFILLER_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1208 U$$934/A1 U$$1218/A2 U$$936/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1209/A sky130_fd_sc_hd__a22o_1
XU$$1219 U$$1219/A U$$1232/A VGND VGND VPWR VPWR U$$1219/X sky130_fd_sc_hd__xor2_1
XFILLER_102_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_81_1 dadda_fa_3_81_1/A dadda_fa_3_81_1/B dadda_fa_3_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/CIN dadda_fa_4_81_2/A sky130_fd_sc_hd__fa_2
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_74_0 dadda_fa_3_74_0/A dadda_fa_3_74_0/B dadda_fa_3_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/B dadda_fa_4_74_1/CIN sky130_fd_sc_hd__fa_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3100 _591_/Q U$$3018/X U$$4335/A1 U$$3019/X VGND VGND VPWR VPWR U$$3101/A sky130_fd_sc_hd__a22o_1
XFILLER_66_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3111 U$$3111/A U$$3137/B VGND VGND VPWR VPWR U$$3111/X sky130_fd_sc_hd__xor2_1
XU$$3122 _602_/Q U$$3018/X _603_/Q U$$3019/X VGND VGND VPWR VPWR U$$3123/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_1 dadda_fa_4_110_1/A dadda_fa_4_110_1/B dadda_fa_4_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/B dadda_fa_5_110_1/B sky130_fd_sc_hd__fa_1
XFILLER_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3133 U$$3133/A U$$3137/B VGND VGND VPWR VPWR U$$3133/X sky130_fd_sc_hd__xor2_1
XU$$3144 U$$4514/A1 U$$3146/A2 U$$4379/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3145/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2410 U$$2410/A U$$2436/B VGND VGND VPWR VPWR U$$2410/X sky130_fd_sc_hd__xor2_1
XU$$3155 U$$3153/Y _662_/Q _661_/Q U$$3154/X U$$3151/Y VGND VGND VPWR VPWR U$$3155/X
+ sky130_fd_sc_hd__a32o_4
Xdadda_fa_2_36_5 input186/X dadda_fa_2_36_5/B dadda_fa_2_36_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_37_2/A dadda_fa_4_36_0/A sky130_fd_sc_hd__fa_2
XU$$2421 U$$914/A1 U$$2421/A2 _595_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2422/A sky130_fd_sc_hd__a22o_1
XU$$3166 U$$3166/A U$$3244/B VGND VGND VPWR VPWR U$$3166/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_0 dadda_fa_4_103_0/A dadda_fa_4_103_0/B dadda_fa_4_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/A dadda_fa_5_103_1/A sky130_fd_sc_hd__fa_1
XU$$3177 _561_/Q U$$3241/A2 U$$28/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3178/A sky130_fd_sc_hd__a22o_1
XU$$2432 U$$2432/A U$$2432/B VGND VGND VPWR VPWR U$$2432/X sky130_fd_sc_hd__xor2_1
XFILLER_62_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2443 U$$799/A1 U$$2463/A2 U$$938/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2444/A sky130_fd_sc_hd__a22o_1
XU$$3188 U$$3188/A U$$3224/B VGND VGND VPWR VPWR U$$3188/X sky130_fd_sc_hd__xor2_1
XU$$2454 U$$2454/A _651_/Q VGND VGND VPWR VPWR U$$2454/X sky130_fd_sc_hd__xor2_1
XU$$1720 U$$2953/A1 U$$1770/A2 _587_/Q U$$1770/B2 VGND VGND VPWR VPWR U$$1721/A sky130_fd_sc_hd__a22o_1
XFILLER_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3199 U$$4156/B1 U$$3241/A2 _573_/Q U$$3253/B2 VGND VGND VPWR VPWR U$$3200/A sky130_fd_sc_hd__a22o_1
XFILLER_50_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2465 _651_/Q VGND VGND VPWR VPWR U$$2465/Y sky130_fd_sc_hd__inv_1
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1731 U$$1731/A U$$1781/A VGND VGND VPWR VPWR U$$1731/X sky130_fd_sc_hd__xor2_1
XU$$2476 U$$8/B1 U$$2574/A2 U$$971/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2477/A sky130_fd_sc_hd__a22o_1
XU$$2487 U$$2487/A U$$2533/B VGND VGND VPWR VPWR U$$2487/X sky130_fd_sc_hd__xor2_1
XU$$1742 U$$98/A1 U$$1648/X U$$98/B1 U$$1649/X VGND VGND VPWR VPWR U$$1743/A sky130_fd_sc_hd__a22o_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1753 U$$1753/A _641_/Q VGND VGND VPWR VPWR U$$1753/X sky130_fd_sc_hd__xor2_1
XU$$2498 U$$30/B1 U$$2534/A2 U$$3457/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2499/A sky130_fd_sc_hd__a22o_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1764 _608_/Q U$$1648/X _609_/Q U$$1649/X VGND VGND VPWR VPWR U$$1765/A sky130_fd_sc_hd__a22o_1
XU$$1775 U$$1775/A U$$1781/A VGND VGND VPWR VPWR U$$1775/X sky130_fd_sc_hd__xor2_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1786 U$$1784/B U$$1781/A _642_/Q U$$1781/Y VGND VGND VPWR VPWR U$$1786/X sky130_fd_sc_hd__a22o_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1797 U$$16/A1 U$$1867/A2 U$$975/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1798/A sky130_fd_sc_hd__a22o_1
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_96_1 dadda_fa_5_96_1/A dadda_fa_5_96_1/B dadda_fa_5_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/B dadda_fa_7_96_0/A sky130_fd_sc_hd__fa_1
XFILLER_174_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput30 a[36] VGND VGND VPWR VPWR _652_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 a[46] VGND VGND VPWR VPWR _662_/D sky130_fd_sc_hd__clkbuf_1
Xinput52 a[56] VGND VGND VPWR VPWR _672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput63 a[8] VGND VGND VPWR VPWR _624_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_128_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_89_0 dadda_fa_5_89_0/A dadda_fa_5_89_0/B dadda_fa_5_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/A dadda_fa_6_89_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_7_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput74 b[18] VGND VGND VPWR VPWR _570_/D sky130_fd_sc_hd__clkbuf_4
Xinput85 b[28] VGND VGND VPWR VPWR _580_/D sky130_fd_sc_hd__clkbuf_4
Xinput96 b[38] VGND VGND VPWR VPWR _590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$405 final_adder.U$$322/B final_adder.U$$630/B final_adder.U$$261/X
+ VGND VGND VPWR VPWR final_adder.U$$634/B sky130_fd_sc_hd__a21o_1
Xrepeater620 U$$4510/A1 VGND VGND VPWR VPWR U$$948/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$427 final_adder.U$$344/B final_adder.U$$718/B final_adder.U$$305/X
+ VGND VGND VPWR VPWR final_adder.U$$722/B sky130_fd_sc_hd__a21o_1
Xrepeater631 _606_/Q VGND VGND VPWR VPWR U$$4500/A1 sky130_fd_sc_hd__buf_12
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater642 _601_/Q VGND VGND VPWR VPWR U$$928/A1 sky130_fd_sc_hd__buf_12
XFILLER_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$449 final_adder.U$$272/B final_adder.U$$654/B final_adder.U$$161/X
+ VGND VGND VPWR VPWR final_adder.U$$656/B sky130_fd_sc_hd__a21o_1
XFILLER_123_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater653 _596_/Q VGND VGND VPWR VPWR U$$96/A1 sky130_fd_sc_hd__buf_12
Xrepeater664 U$$908/A1 VGND VGND VPWR VPWR U$$86/A1 sky130_fd_sc_hd__buf_12
Xrepeater675 _587_/Q VGND VGND VPWR VPWR U$$78/A1 sky130_fd_sc_hd__buf_12
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater686 U$$892/A1 VGND VGND VPWR VPWR U$$68/B1 sky130_fd_sc_hd__buf_12
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater697 U$$4446/A1 VGND VGND VPWR VPWR U$$3624/A1 sky130_fd_sc_hd__buf_12
XU$$4390 U$$4390/A1 U$$4388/X _552_/Q U$$4389/X VGND VGND VPWR VPWR U$$4391/A sky130_fd_sc_hd__a22o_1
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_91_0 dadda_fa_4_91_0/A dadda_fa_4_91_0/B dadda_fa_4_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/A dadda_fa_5_91_1/A sky130_fd_sc_hd__fa_1
XFILLER_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_105_2 U$$4473/X input135/X dadda_fa_3_105_2/CIN VGND VGND VPWR VPWR dadda_fa_4_106_1/A
+ dadda_fa_4_105_2/B sky130_fd_sc_hd__fa_1
XFILLER_161_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_789__841 VGND VGND VPWR VPWR _789__841/HI U$$4423/B sky130_fd_sc_hd__conb_1
XFILLER_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_119_0 dadda_fa_6_119_0/A dadda_fa_6_119_0/B dadda_fa_6_119_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_120_0/B dadda_fa_7_119_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$800 U$$800/A U$$822/A VGND VGND VPWR VPWR U$$800/X sky130_fd_sc_hd__xor2_1
X_673_ _677_/CLK _673_/D VGND VGND VPWR VPWR _673_/Q sky130_fd_sc_hd__dfxtp_4
XU$$811 U$$948/A1 U$$817/A2 U$$950/A1 U$$817/B2 VGND VGND VPWR VPWR U$$812/A sky130_fd_sc_hd__a22o_1
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$822 U$$822/A VGND VGND VPWR VPWR U$$822/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_3_39_3 dadda_fa_3_39_3/A dadda_fa_3_39_3/B dadda_fa_3_39_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/B dadda_fa_4_39_2/CIN sky130_fd_sc_hd__fa_2
XU$$833 U$$833/A U$$923/B VGND VGND VPWR VPWR U$$833/X sky130_fd_sc_hd__xor2_1
XU$$844 _559_/Q U$$910/A2 U$$983/A1 U$$910/B2 VGND VGND VPWR VPWR U$$845/A sky130_fd_sc_hd__a22o_1
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$855 U$$855/A U$$903/B VGND VGND VPWR VPWR U$$855/X sky130_fd_sc_hd__xor2_1
XU$$866 _570_/Q U$$928/A2 U$$46/A1 U$$928/B2 VGND VGND VPWR VPWR U$$867/A sky130_fd_sc_hd__a22o_1
XU$$1005 U$$868/A1 U$$999/A2 U$$48/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1006/A sky130_fd_sc_hd__a22o_1
XU$$1016 U$$1016/A U$$980/B VGND VGND VPWR VPWR U$$1016/X sky130_fd_sc_hd__xor2_1
XU$$877 U$$877/A U$$943/B VGND VGND VPWR VPWR U$$877/X sky130_fd_sc_hd__xor2_1
XU$$888 U$$66/A1 U$$910/A2 U$$68/A1 U$$910/B2 VGND VGND VPWR VPWR U$$889/A sky130_fd_sc_hd__a22o_1
XFILLER_73_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1027 U$$68/A1 U$$999/A2 U$$68/B1 U$$987/B2 VGND VGND VPWR VPWR U$$1028/A sky130_fd_sc_hd__a22o_1
XU$$1038 U$$1038/A U$$998/B VGND VGND VPWR VPWR U$$1038/X sky130_fd_sc_hd__xor2_1
XU$$899 U$$899/A U$$903/B VGND VGND VPWR VPWR U$$899/X sky130_fd_sc_hd__xor2_1
XFILLER_71_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1049 U$$912/A1 U$$1093/A2 U$$914/A1 U$$1073/B2 VGND VGND VPWR VPWR U$$1050/A sky130_fd_sc_hd__a22o_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_28_3 U$$1260/X U$$1393/X VGND VGND VPWR VPWR dadda_fa_3_29_2/CIN dadda_fa_4_28_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_41_3 U$$2749/X input192/X dadda_fa_2_41_3/CIN VGND VGND VPWR VPWR dadda_fa_3_42_1/B
+ dadda_fa_3_41_3/B sky130_fd_sc_hd__fa_2
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_34_2 U$$1139/X U$$1272/X U$$1405/X VGND VGND VPWR VPWR dadda_fa_3_35_1/A
+ dadda_fa_3_34_3/A sky130_fd_sc_hd__fa_1
XU$$2240 U$$48/A1 U$$2270/A2 U$$50/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2241/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_1 dadda_fa_5_11_1/A dadda_fa_5_11_1/B dadda_ha_4_11_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_12_0/B dadda_fa_7_11_0/A sky130_fd_sc_hd__fa_2
XU$$2251 U$$2251/A U$$2257/B VGND VGND VPWR VPWR U$$2251/X sky130_fd_sc_hd__xor2_1
XU$$2262 U$$70/A1 U$$2196/X U$$70/B1 U$$2197/X VGND VGND VPWR VPWR U$$2263/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_27_1 U$$460/X U$$593/X U$$726/X VGND VGND VPWR VPWR dadda_fa_3_28_2/B
+ dadda_fa_3_27_3/CIN sky130_fd_sc_hd__fa_1
XU$$2273 U$$2273/A U$$2327/B VGND VGND VPWR VPWR U$$2273/X sky130_fd_sc_hd__xor2_1
XFILLER_90_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2284 U$$914/A1 U$$2316/A2 U$$92/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2285/A sky130_fd_sc_hd__a22o_1
XU$$2295 U$$2295/A _649_/Q VGND VGND VPWR VPWR U$$2295/X sky130_fd_sc_hd__xor2_1
XU$$1550 U$$1550/A U$$1580/B VGND VGND VPWR VPWR U$$1550/X sky130_fd_sc_hd__xor2_1
XU$$1561 U$$876/A1 U$$1591/A2 U$$878/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1562/A sky130_fd_sc_hd__a22o_1
XFILLER_22_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1572 U$$1572/A U$$1643/A VGND VGND VPWR VPWR U$$1572/X sky130_fd_sc_hd__xor2_1
XU$$1583 U$$2953/A1 U$$1605/A2 U$$76/B1 U$$1605/B2 VGND VGND VPWR VPWR U$$1584/A sky130_fd_sc_hd__a22o_1
XU$$1594 U$$1594/A U$$1614/B VGND VGND VPWR VPWR U$$1594/X sky130_fd_sc_hd__xor2_1
XFILLER_187_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_79_4 U$$2692/X U$$2825/X U$$2958/X VGND VGND VPWR VPWR dadda_fa_2_80_1/CIN
+ dadda_fa_2_79_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$202 final_adder.U$$697/A final_adder.U$$696/A VGND VGND VPWR VPWR
+ final_adder.U$$292/A sky130_fd_sc_hd__and2_1
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$213 final_adder.U$$707/A final_adder.U$$579/B1 final_adder.U$$213/B1
+ VGND VGND VPWR VPWR final_adder.U$$213/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$224 final_adder.U$$719/A final_adder.U$$718/A VGND VGND VPWR VPWR
+ final_adder.U$$304/B sky130_fd_sc_hd__and2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_2 dadda_fa_4_49_2/A dadda_fa_4_49_2/B dadda_fa_4_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/CIN dadda_fa_5_49_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$235 final_adder.U$$729/A final_adder.U$$601/B1 final_adder.U$$235/B1
+ VGND VGND VPWR VPWR final_adder.U$$235/X sky130_fd_sc_hd__a21o_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$246 final_adder.U$$741/A final_adder.U$$740/A VGND VGND VPWR VPWR
+ final_adder.U$$314/A sky130_fd_sc_hd__and2_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater450 U$$1100/X VGND VGND VPWR VPWR U$$1200/A2 sky130_fd_sc_hd__buf_12
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$257 final_adder.U$$130/X final_adder.U$$624/B final_adder.U$$131/X
+ VGND VGND VPWR VPWR final_adder.U$$626/B sky130_fd_sc_hd__a21o_2
Xrepeater461 U$$4115/X VGND VGND VPWR VPWR U$$4244/B2 sky130_fd_sc_hd__buf_12
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$268 final_adder.U$$268/A final_adder.U$$268/B VGND VGND VPWR VPWR
+ final_adder.U$$326/B sky130_fd_sc_hd__and2_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$107 U$$107/A U$$89/B VGND VGND VPWR VPWR U$$107/X sky130_fd_sc_hd__xor2_1
Xrepeater472 U$$3545/B2 VGND VGND VPWR VPWR U$$3525/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$279 final_adder.U$$278/A final_adder.U$$173/X final_adder.U$$175/X
+ VGND VGND VPWR VPWR final_adder.U$$279/X sky130_fd_sc_hd__a21o_1
XU$$118 U$$940/A1 U$$4/X U$$942/A1 U$$5/X VGND VGND VPWR VPWR U$$119/A sky130_fd_sc_hd__a22o_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater483 U$$2745/X VGND VGND VPWR VPWR U$$2826/B2 sky130_fd_sc_hd__buf_12
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_19_0 dadda_fa_7_19_0/A dadda_fa_7_19_0/B dadda_fa_7_19_0/CIN VGND VGND
+ VPWR VPWR _444_/D _315_/D sky130_fd_sc_hd__fa_2
XU$$129 U$$129/A _617_/Q VGND VGND VPWR VPWR U$$129/X sky130_fd_sc_hd__xor2_1
Xrepeater494 U$$2060/X VGND VGND VPWR VPWR U$$2117/B2 sky130_fd_sc_hd__buf_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_110_0 _698__918/HI U$$3286/X U$$3419/X VGND VGND VPWR VPWR dadda_fa_4_111_0/CIN
+ dadda_fa_4_110_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput220 c[67] VGND VGND VPWR VPWR input220/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput231 c[77] VGND VGND VPWR VPWR input231/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput242 c[87] VGND VGND VPWR VPWR input242/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_51_2 dadda_fa_3_51_2/A dadda_fa_3_51_2/B dadda_fa_3_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/A dadda_fa_4_51_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_67_2 U$$939/X U$$1072/X U$$1205/X VGND VGND VPWR VPWR dadda_fa_1_68_6/A
+ dadda_fa_1_67_8/A sky130_fd_sc_hd__fa_1
Xinput253 c[97] VGND VGND VPWR VPWR input253/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_44_1 dadda_fa_3_44_1/A dadda_fa_3_44_1/B dadda_fa_3_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/CIN dadda_fa_4_44_2/A sky130_fd_sc_hd__fa_2
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_21_0 dadda_fa_6_21_0/A dadda_fa_6_21_0/B dadda_fa_6_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_22_0/B dadda_fa_7_21_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_37_0 dadda_fa_3_37_0/A dadda_fa_3_37_0/B dadda_fa_3_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/B dadda_fa_4_37_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_656_ _656_/CLK _656_/D VGND VGND VPWR VPWR _656_/Q sky130_fd_sc_hd__dfxtp_1
XU$$630 U$$630/A1 U$$682/A2 U$$84/A1 U$$553/X VGND VGND VPWR VPWR U$$631/A sky130_fd_sc_hd__a22o_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$641 U$$641/A U$$661/B VGND VGND VPWR VPWR U$$641/X sky130_fd_sc_hd__xor2_1
XFILLER_16_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$652 U$$926/A1 U$$682/A2 U$$928/A1 U$$553/X VGND VGND VPWR VPWR U$$653/A sky130_fd_sc_hd__a22o_1
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$663 U$$663/A _625_/Q VGND VGND VPWR VPWR U$$663/X sky130_fd_sc_hd__xor2_1
XFILLER_189_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$674 U$$948/A1 U$$682/A2 U$$950/A1 U$$553/X VGND VGND VPWR VPWR U$$675/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$685 _625_/Q VGND VGND VPWR VPWR U$$685/Y sky130_fd_sc_hd__inv_1
XFILLER_72_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_587_ _594_/CLK _587_/D VGND VGND VPWR VPWR _587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$696 U$$696/A U$$778/B VGND VGND VPWR VPWR U$$696/X sky130_fd_sc_hd__xor2_1
XFILLER_189_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_96_4 U$$4056/X U$$4189/X U$$4322/X VGND VGND VPWR VPWR dadda_fa_3_97_1/CIN
+ dadda_fa_3_96_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_89_3 input244/X dadda_fa_2_89_3/B dadda_fa_2_89_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_90_1/B dadda_fa_3_89_3/B sky130_fd_sc_hd__fa_2
XFILLER_141_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_59_1 dadda_fa_5_59_1/A dadda_fa_5_59_1/B dadda_fa_5_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/B dadda_fa_7_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_113_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_105_1 U$$3276/X U$$3409/X U$$3542/X VGND VGND VPWR VPWR dadda_fa_3_106_3/B
+ dadda_fa_4_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2070 U$$2070/A U$$2118/B VGND VGND VPWR VPWR U$$2070/X sky130_fd_sc_hd__xor2_1
XU$$2081 U$$26/A1 U$$2117/A2 U$$987/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2082/A sky130_fd_sc_hd__a22o_1
XU$$2092 U$$2092/A U$$2118/B VGND VGND VPWR VPWR U$$2092/X sky130_fd_sc_hd__xor2_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1380 U$$8/B1 U$$1474/A2 U$$971/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1381/A sky130_fd_sc_hd__a22o_1
XU$$1391 U$$1391/A U$$1479/B VGND VGND VPWR VPWR U$$1391/X sky130_fd_sc_hd__xor2_1
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_84_2 U$$2170/X U$$2303/X U$$2436/X VGND VGND VPWR VPWR dadda_fa_2_85_2/CIN
+ dadda_fa_2_84_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_61_1 dadda_fa_4_61_1/A dadda_fa_4_61_1/B dadda_fa_4_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/B dadda_fa_5_61_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_1 U$$1757/X U$$1890/X U$$2023/X VGND VGND VPWR VPWR dadda_fa_2_78_0/CIN
+ dadda_fa_2_77_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_54_0 dadda_fa_4_54_0/A dadda_fa_4_54_0/B dadda_fa_4_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/A dadda_fa_5_54_1/A sky130_fd_sc_hd__fa_1
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_510_ _510_/CLK _510_/D VGND VGND VPWR VPWR _510_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ _461_/CLK _441_/D VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _501_/CLK _372_/D VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_99_2 dadda_fa_3_99_2/A dadda_fa_3_99_2/B dadda_fa_3_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/A dadda_fa_4_99_2/B sky130_fd_sc_hd__fa_1
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_69_0 dadda_fa_6_69_0/A dadda_fa_6_69_0/B dadda_fa_6_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_70_0/B dadda_fa_7_69_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_72_0 _682__902/HI U$$683/X U$$816/X VGND VGND VPWR VPWR dadda_fa_1_73_7/A
+ dadda_fa_1_72_8/A sky130_fd_sc_hd__fa_1
XFILLER_122_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$460 U$$460/A U$$530/B VGND VGND VPWR VPWR U$$460/X sky130_fd_sc_hd__xor2_2
X_639_ _639_/CLK _639_/D VGND VGND VPWR VPWR _639_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$471 U$$60/A1 U$$491/A2 U$$62/A1 U$$416/X VGND VGND VPWR VPWR U$$472/A sky130_fd_sc_hd__a22o_1
XU$$482 U$$482/A _623_/Q VGND VGND VPWR VPWR U$$482/X sky130_fd_sc_hd__xor2_1
XFILLER_189_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$493 U$$82/A1 U$$545/A2 U$$84/A1 U$$416/X VGND VGND VPWR VPWR U$$494/A sky130_fd_sc_hd__a22o_1
XFILLER_60_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_94_1 U$$3121/X U$$3254/X U$$3387/X VGND VGND VPWR VPWR dadda_fa_3_95_0/CIN
+ dadda_fa_3_94_2/CIN sky130_fd_sc_hd__fa_1
X_735__787 VGND VGND VPWR VPWR _735__787/HI U$$2600/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_5_71_0 dadda_fa_5_71_0/A dadda_fa_5_71_0/B dadda_fa_5_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/A dadda_fa_6_71_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_87_0 U$$3639/X U$$3772/X U$$3905/X VGND VGND VPWR VPWR dadda_fa_3_88_0/B
+ dadda_fa_3_87_2/B sky130_fd_sc_hd__fa_1
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_70_8 dadda_fa_1_70_8/A dadda_fa_1_70_8/B dadda_fa_1_70_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_3/A dadda_fa_3_70_0/A sky130_fd_sc_hd__fa_2
XFILLER_86_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_63_7 dadda_fa_1_63_7/A dadda_fa_1_63_7/B dadda_fa_1_63_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/CIN dadda_fa_2_63_5/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_6 U$$3577/X U$$3710/X U$$3843/X VGND VGND VPWR VPWR dadda_fa_2_57_2/B
+ dadda_fa_2_56_5/B sky130_fd_sc_hd__fa_1
XFILLER_67_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_49_5 U$$2100/X U$$2233/X U$$2366/X VGND VGND VPWR VPWR dadda_fa_2_50_2/B
+ dadda_fa_2_49_5/B sky130_fd_sc_hd__fa_2
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_8_0 dadda_fa_7_8_0/A dadda_fa_7_8_0/B dadda_fa_7_8_0/CIN VGND VGND VPWR
+ VPWR _433_/D _304_/D sky130_fd_sc_hd__fa_2
XFILLER_39_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_86_0 dadda_fa_7_86_0/A dadda_fa_7_86_0/B dadda_fa_7_86_0/CIN VGND VGND
+ VPWR VPWR _511_/D _382_/D sky130_fd_sc_hd__fa_1
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_684__904 VGND VGND VPWR VPWR _684__904/HI _684__904/LO sky130_fd_sc_hd__conb_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4208 U$$98/A1 U$$4244/A2 U$$4484/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4209/A sky130_fd_sc_hd__a22o_1
XU$$4219 U$$4219/A U$$4246/A VGND VGND VPWR VPWR U$$4219/X sky130_fd_sc_hd__xor2_1
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3507 _589_/Q U$$3545/A2 _590_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3508/A sky130_fd_sc_hd__a22o_1
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3518 U$$3518/A _667_/Q VGND VGND VPWR VPWR U$$3518/X sky130_fd_sc_hd__xor2_1
XFILLER_86_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_101_0 dadda_fa_6_101_0/A dadda_fa_6_101_0/B dadda_fa_6_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_102_0/B dadda_fa_7_101_0/CIN sky130_fd_sc_hd__fa_1
XU$$3529 _600_/Q U$$3545/A2 _601_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3530/A sky130_fd_sc_hd__a22o_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2806 U$$3489/B1 U$$2870/A2 U$$4178/A1 U$$2834/B2 VGND VGND VPWR VPWR U$$2807/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2817 U$$2817/A U$$2839/B VGND VGND VPWR VPWR U$$2817/X sky130_fd_sc_hd__xor2_1
XFILLER_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2828 U$$4335/A1 U$$2868/A2 _593_/Q U$$2870/B2 VGND VGND VPWR VPWR U$$2829/A sky130_fd_sc_hd__a22o_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2839 U$$2839/A U$$2839/B VGND VGND VPWR VPWR U$$2839/X sky130_fd_sc_hd__xor2_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_424_ _447_/CLK _424_/D VGND VGND VPWR VPWR _424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_355_ _490_/CLK _355_/D VGND VGND VPWR VPWR _355_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_286_ _612_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_66_5 dadda_fa_2_66_5/A dadda_fa_2_66_5/B dadda_fa_2_66_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_2/A dadda_fa_4_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_59_4 dadda_fa_2_59_4/A dadda_fa_2_59_4/B dadda_fa_2_59_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/CIN dadda_fa_3_59_3/CIN sky130_fd_sc_hd__fa_2
Xinput6 a[14] VGND VGND VPWR VPWR _630_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$290 U$$16/A1 U$$278/X U$$975/B1 U$$279/X VGND VGND VPWR VPWR U$$291/A sky130_fd_sc_hd__a22o_1
XFILLER_189_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$4 _428_/Q _300_/Q VGND VGND VPWR VPWR final_adder.U$$499/B1 final_adder.U$$626/A
+ sky130_fd_sc_hd__ha_2
XFILLER_133_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput310 _200_/Q VGND VGND VPWR VPWR o[32] sky130_fd_sc_hd__buf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 _210_/Q VGND VGND VPWR VPWR o[42] sky130_fd_sc_hd__buf_2
Xoutput332 _220_/Q VGND VGND VPWR VPWR o[52] sky130_fd_sc_hd__buf_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 _230_/Q VGND VGND VPWR VPWR o[62] sky130_fd_sc_hd__buf_2
Xoutput354 _240_/Q VGND VGND VPWR VPWR o[72] sky130_fd_sc_hd__buf_2
Xoutput365 _250_/Q VGND VGND VPWR VPWR o[82] sky130_fd_sc_hd__buf_2
Xoutput376 _260_/Q VGND VGND VPWR VPWR o[92] sky130_fd_sc_hd__buf_2
XFILLER_114_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_61_4 U$$3587/X U$$3720/X U$$3853/X VGND VGND VPWR VPWR dadda_fa_2_62_1/CIN
+ dadda_fa_2_61_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_709__929 VGND VGND VPWR VPWR _709__929/HI _709__929/LO sky130_fd_sc_hd__conb_1
XFILLER_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_54_3 U$$1977/X U$$2110/X U$$2243/X VGND VGND VPWR VPWR dadda_fa_2_55_1/B
+ dadda_fa_2_54_4/B sky130_fd_sc_hd__fa_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_31_2 dadda_fa_4_31_2/A dadda_fa_4_31_2/B dadda_fa_4_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/CIN dadda_fa_5_31_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_47_2 U$$899/X U$$1032/X U$$1165/X VGND VGND VPWR VPWR dadda_fa_2_48_2/A
+ dadda_fa_2_47_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_24_1 dadda_fa_4_24_1/A dadda_fa_4_24_1/B dadda_fa_4_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/B dadda_fa_5_24_1/B sky130_fd_sc_hd__fa_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_0 U$$706/X U$$839/X U$$972/X VGND VGND VPWR VPWR dadda_fa_5_18_0/A
+ dadda_fa_5_17_1/A sky130_fd_sc_hd__fa_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_69_3 dadda_fa_3_69_3/A dadda_fa_3_69_3/B dadda_fa_3_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/B dadda_fa_4_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4005 _564_/Q U$$3977/X _565_/Q U$$3978/X VGND VGND VPWR VPWR U$$4006/A sky130_fd_sc_hd__a22o_1
XU$$4016 U$$4016/A U$$4109/A VGND VGND VPWR VPWR U$$4016/X sky130_fd_sc_hd__xor2_1
XU$$4027 _575_/Q U$$4045/A2 U$$4303/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$4028/A sky130_fd_sc_hd__a22o_1
XFILLER_24_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4038 U$$4038/A _675_/Q VGND VGND VPWR VPWR U$$4038/X sky130_fd_sc_hd__xor2_1
XU$$3304 _556_/Q U$$3396/A2 U$$4265/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3305/A sky130_fd_sc_hd__a22o_1
XU$$4049 U$$759/B1 U$$4107/A2 U$$78/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4050/A sky130_fd_sc_hd__a22o_1
XU$$3315 U$$3315/A U$$3397/B VGND VGND VPWR VPWR U$$3315/X sky130_fd_sc_hd__xor2_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3326 _567_/Q U$$3412/A2 U$$40/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3327/A sky130_fd_sc_hd__a22o_1
XU$$3337 U$$3337/A U$$3397/B VGND VGND VPWR VPWR U$$3337/X sky130_fd_sc_hd__xor2_1
XU$$2603 U$$2603/A VGND VGND VPWR VPWR U$$2603/Y sky130_fd_sc_hd__inv_1
XFILLER_74_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3348 U$$4170/A1 U$$3396/A2 U$$3624/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3349/A
+ sky130_fd_sc_hd__a22o_1
XU$$2614 U$$2614/A U$$2710/B VGND VGND VPWR VPWR U$$2614/X sky130_fd_sc_hd__xor2_1
XU$$3359 U$$3359/A U$$3397/B VGND VGND VPWR VPWR U$$3359/X sky130_fd_sc_hd__xor2_1
XU$$2625 U$$979/B1 U$$2667/A2 U$$4271/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2626/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2636 U$$2636/A U$$2694/B VGND VGND VPWR VPWR U$$2636/X sky130_fd_sc_hd__xor2_1
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2647 U$$4289/B1 U$$2607/X U$$4291/B1 U$$2608/X VGND VGND VPWR VPWR U$$2648/A sky130_fd_sc_hd__a22o_1
XU$$1902 U$$1902/A U$$1904/B VGND VGND VPWR VPWR U$$1902/X sky130_fd_sc_hd__xor2_1
XFILLER_34_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1913 U$$952/B1 U$$1785/X U$$956/A1 U$$1786/X VGND VGND VPWR VPWR U$$1914/A sky130_fd_sc_hd__a22o_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2658 U$$2658/A U$$2694/B VGND VGND VPWR VPWR U$$2658/X sky130_fd_sc_hd__xor2_1
XU$$1924 U$$1924/A1 U$$1922/X U$$8/A1 U$$1923/X VGND VGND VPWR VPWR U$$1925/A sky130_fd_sc_hd__a22o_1
XFILLER_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2669 U$$3489/B1 U$$2729/A2 U$$3217/B1 U$$2729/B2 VGND VGND VPWR VPWR U$$2670/A
+ sky130_fd_sc_hd__a22o_1
XU$$1935 U$$1935/A U$$1991/B VGND VGND VPWR VPWR U$$1935/X sky130_fd_sc_hd__xor2_1
XU$$1946 U$$28/A1 U$$1922/X U$$28/B1 U$$1923/X VGND VGND VPWR VPWR U$$1947/A sky130_fd_sc_hd__a22o_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1957 U$$1957/A U$$1991/B VGND VGND VPWR VPWR U$$1957/X sky130_fd_sc_hd__xor2_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1968 U$$735/A1 U$$1922/X U$$52/A1 U$$1923/X VGND VGND VPWR VPWR U$$1969/A sky130_fd_sc_hd__a22o_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _535_/CLK _407_/D VGND VGND VPWR VPWR _407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1979 U$$1979/A U$$1991/B VGND VGND VPWR VPWR U$$1979/X sky130_fd_sc_hd__xor2_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ _469_/CLK _338_/D VGND VGND VPWR VPWR _338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_269_ _280_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_71_3 dadda_fa_2_71_3/A dadda_fa_2_71_3/B dadda_fa_2_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/B dadda_fa_3_71_3/B sky130_fd_sc_hd__fa_1
XFILLER_123_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_64_2 dadda_fa_2_64_2/A dadda_fa_2_64_2/B dadda_fa_2_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/A dadda_fa_3_64_3/A sky130_fd_sc_hd__fa_1
XFILLER_97_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$609 final_adder.U$$736/A final_adder.U$$736/B final_adder.U$$609/B1
+ VGND VGND VPWR VPWR final_adder.U$$737/B sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_41_1 dadda_fa_5_41_1/A dadda_fa_5_41_1/B dadda_fa_5_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/B dadda_fa_7_41_0/A sky130_fd_sc_hd__fa_2
X_847__899 VGND VGND VPWR VPWR _847__899/HI _847__899/LO sky130_fd_sc_hd__conb_1
Xdadda_fa_2_57_1 dadda_fa_2_57_1/A dadda_fa_2_57_1/B dadda_fa_2_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/CIN dadda_fa_3_57_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_34_0 dadda_fa_5_34_0/A dadda_fa_5_34_0/B dadda_fa_5_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/A dadda_fa_6_34_0/CIN sky130_fd_sc_hd__fa_1
XU$$20 U$$20/A1 U$$4/X _559_/Q U$$5/X VGND VGND VPWR VPWR U$$21/A sky130_fd_sc_hd__a22o_1
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$31 U$$31/A U$$9/B VGND VGND VPWR VPWR U$$31/X sky130_fd_sc_hd__xor2_1
XU$$42 _569_/Q U$$4/X _570_/Q U$$5/X VGND VGND VPWR VPWR U$$43/A sky130_fd_sc_hd__a22o_1
XU$$53 U$$53/A U$$3/A VGND VGND VPWR VPWR U$$53/X sky130_fd_sc_hd__xor2_1
XFILLER_38_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$64 U$$64/A1 U$$4/X U$$66/A1 U$$5/X VGND VGND VPWR VPWR U$$65/A sky130_fd_sc_hd__a22o_1
XU$$3860 _560_/Q U$$3912/A2 _561_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3861/A sky130_fd_sc_hd__a22o_1
XU$$75 U$$75/A U$$9/B VGND VGND VPWR VPWR U$$75/X sky130_fd_sc_hd__xor2_1
XU$$3871 U$$3871/A U$$3929/B VGND VGND VPWR VPWR U$$3871/X sky130_fd_sc_hd__xor2_1
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$86 U$$86/A1 U$$4/X U$$88/A1 U$$5/X VGND VGND VPWR VPWR U$$87/A sky130_fd_sc_hd__a22o_1
XU$$3882 _571_/Q U$$3970/A2 _572_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3883/A sky130_fd_sc_hd__a22o_1
XU$$97 U$$97/A U$$3/A VGND VGND VPWR VPWR U$$97/X sky130_fd_sc_hd__xor2_1
XFILLER_53_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3893 U$$3893/A U$$3893/B VGND VGND VPWR VPWR U$$3893/X sky130_fd_sc_hd__xor2_1
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_750__802 VGND VGND VPWR VPWR _750__802/HI U$$3431/A1 sky130_fd_sc_hd__conb_1
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_79_2 dadda_fa_4_79_2/A dadda_fa_4_79_2/B dadda_fa_4_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/CIN dadda_fa_5_79_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_49_0 dadda_fa_7_49_0/A dadda_fa_7_49_0/B dadda_fa_7_49_0/CIN VGND VGND
+ VPWR VPWR _474_/D _345_/D sky130_fd_sc_hd__fa_2
XFILLER_48_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_52_0 U$$377/X U$$510/X U$$643/X VGND VGND VPWR VPWR dadda_fa_2_53_0/B
+ dadda_fa_2_52_3/B sky130_fd_sc_hd__fa_2
XFILLER_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1209 U$$1209/A _633_/Q VGND VGND VPWR VPWR U$$1209/X sky130_fd_sc_hd__xor2_1
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_50_clk _536_/CLK VGND VGND VPWR VPWR _601_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_81_2 dadda_fa_3_81_2/A dadda_fa_3_81_2/B dadda_fa_3_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/A dadda_fa_4_81_2/B sky130_fd_sc_hd__fa_1
XFILLER_139_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_74_1 dadda_fa_3_74_1/A dadda_fa_3_74_1/B dadda_fa_3_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/CIN dadda_fa_4_74_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_51_0 dadda_fa_6_51_0/A dadda_fa_6_51_0/B dadda_fa_6_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_52_0/B dadda_fa_7_51_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_67_0 dadda_fa_3_67_0/A dadda_fa_3_67_0/B dadda_fa_3_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/B dadda_fa_4_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3101 U$$3101/A U$$3137/B VGND VGND VPWR VPWR U$$3101/X sky130_fd_sc_hd__xor2_1
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3112 U$$96/B1 U$$3018/X U$$785/A1 U$$3019/X VGND VGND VPWR VPWR U$$3113/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_2 dadda_fa_4_110_2/A dadda_fa_4_110_2/B dadda_ha_3_110_3/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/CIN dadda_fa_5_110_1/CIN sky130_fd_sc_hd__fa_1
XU$$3123 U$$3123/A U$$3137/B VGND VGND VPWR VPWR U$$3123/X sky130_fd_sc_hd__xor2_1
XU$$3134 U$$4504/A1 U$$3018/X U$$4506/A1 U$$3019/X VGND VGND VPWR VPWR U$$3135/A sky130_fd_sc_hd__a22o_1
XU$$2400 U$$2400/A U$$2464/B VGND VGND VPWR VPWR U$$2400/X sky130_fd_sc_hd__xor2_1
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3145 U$$3145/A _661_/Q VGND VGND VPWR VPWR U$$3145/X sky130_fd_sc_hd__xor2_1
XU$$2411 _589_/Q U$$2421/A2 _590_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2412/A sky130_fd_sc_hd__a22o_1
XFILLER_19_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3156 U$$3154/B _661_/Q _662_/Q U$$3151/Y VGND VGND VPWR VPWR U$$3156/X sky130_fd_sc_hd__a22o_4
XU$$2422 U$$2422/A U$$2436/B VGND VGND VPWR VPWR U$$2422/X sky130_fd_sc_hd__xor2_1
XFILLER_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_103_1 dadda_fa_4_103_1/A dadda_fa_4_103_1/B dadda_fa_4_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/B dadda_fa_5_103_1/B sky130_fd_sc_hd__fa_1
XU$$3167 _556_/Q U$$3243/A2 U$$4265/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3168/A sky130_fd_sc_hd__a22o_1
XU$$2433 _600_/Q U$$2463/A2 U$$928/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2434/A sky130_fd_sc_hd__a22o_1
XU$$3178 U$$3178/A U$$3224/B VGND VGND VPWR VPWR U$$3178/X sky130_fd_sc_hd__xor2_1
XU$$2444 U$$2444/A U$$2464/B VGND VGND VPWR VPWR U$$2444/X sky130_fd_sc_hd__xor2_1
XU$$3189 U$$4285/A1 U$$3241/A2 U$$3191/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3190/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1710 U$$3489/B1 U$$1726/A2 U$$3217/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1711/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2455 U$$4510/A1 U$$2463/A2 U$$950/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2456/A
+ sky130_fd_sc_hd__a22o_1
XU$$1721 U$$1721/A _641_/Q VGND VGND VPWR VPWR U$$1721/X sky130_fd_sc_hd__xor2_1
XU$$2466 _651_/Q VGND VGND VPWR VPWR U$$2466/Y sky130_fd_sc_hd__inv_1
XU$$1732 U$$771/B1 U$$1734/A2 U$$90/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1733/A sky130_fd_sc_hd__a22o_1
XU$$2477 U$$2477/A U$$2533/B VGND VGND VPWR VPWR U$$2477/X sky130_fd_sc_hd__xor2_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1743 U$$1743/A U$$1781/A VGND VGND VPWR VPWR U$$1743/X sky130_fd_sc_hd__xor2_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2488 U$$979/B1 U$$2534/A2 U$$4271/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2489/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1754 U$$932/A1 U$$1648/X U$$934/A1 U$$1649/X VGND VGND VPWR VPWR U$$1755/A sky130_fd_sc_hd__a22o_1
XU$$2499 U$$2499/A U$$2533/B VGND VGND VPWR VPWR U$$2499/X sky130_fd_sc_hd__xor2_1
XU$$1765 U$$1765/A _641_/Q VGND VGND VPWR VPWR U$$1765/X sky130_fd_sc_hd__xor2_1
XFILLER_159_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1776 U$$4379/A1 U$$1648/X U$$956/A1 U$$1649/X VGND VGND VPWR VPWR U$$1777/A sky130_fd_sc_hd__a22o_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1787 U$$1787/A1 U$$1867/A2 U$$8/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1788/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_124_0 dadda_fa_7_124_0/A dadda_fa_7_124_0/B dadda_fa_7_124_0/CIN VGND
+ VGND VPWR VPWR _549_/D _420_/D sky130_fd_sc_hd__fa_2
XU$$1798 U$$1798/A U$$1918/A VGND VGND VPWR VPWR U$$1798/X sky130_fd_sc_hd__xor2_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_187_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 a[27] VGND VGND VPWR VPWR _643_/D sky130_fd_sc_hd__clkbuf_4
Xinput31 a[37] VGND VGND VPWR VPWR _653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 a[47] VGND VGND VPWR VPWR _663_/D sky130_fd_sc_hd__clkbuf_1
Xinput53 a[57] VGND VGND VPWR VPWR _673_/D sky130_fd_sc_hd__clkbuf_1
Xinput64 a[9] VGND VGND VPWR VPWR _625_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_156_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_89_1 dadda_fa_5_89_1/A dadda_fa_5_89_1/B dadda_fa_5_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/B dadda_fa_7_89_0/A sky130_fd_sc_hd__fa_1
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput75 b[19] VGND VGND VPWR VPWR _571_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput86 b[29] VGND VGND VPWR VPWR _581_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_143_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 b[39] VGND VGND VPWR VPWR _591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater610 _617_/Q VGND VGND VPWR VPWR U$$3/A sky130_fd_sc_hd__buf_12
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$417 final_adder.U$$334/B final_adder.U$$678/B final_adder.U$$285/X
+ VGND VGND VPWR VPWR final_adder.U$$682/B sky130_fd_sc_hd__a21o_1
Xrepeater621 _611_/Q VGND VGND VPWR VPWR U$$4510/A1 sky130_fd_sc_hd__buf_12
XFILLER_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater632 _605_/Q VGND VGND VPWR VPWR U$$936/A1 sky130_fd_sc_hd__buf_12
Xrepeater643 _600_/Q VGND VGND VPWR VPWR U$$926/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$439 final_adder.U$$262/B final_adder.U$$634/B final_adder.U$$141/X
+ VGND VGND VPWR VPWR final_adder.U$$636/B sky130_fd_sc_hd__a21o_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater654 _595_/Q VGND VGND VPWR VPWR U$$92/B1 sky130_fd_sc_hd__buf_12
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater665 U$$908/A1 VGND VGND VPWR VPWR U$$771/A1 sky130_fd_sc_hd__buf_12
Xrepeater676 _587_/Q VGND VGND VPWR VPWR U$$76/B1 sky130_fd_sc_hd__buf_12
XFILLER_26_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater687 U$$70/A1 VGND VGND VPWR VPWR U$$892/A1 sky130_fd_sc_hd__buf_12
XFILLER_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4380 U$$4380/A _679_/Q VGND VGND VPWR VPWR U$$4380/X sky130_fd_sc_hd__xor2_2
Xrepeater698 _579_/Q VGND VGND VPWR VPWR U$$4446/A1 sky130_fd_sc_hd__buf_12
XU$$4391 U$$4391/A U$$4391/B VGND VGND VPWR VPWR U$$4391/X sky130_fd_sc_hd__xor2_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3690 U$$539/A1 U$$3566/X _613_/Q U$$3567/X VGND VGND VPWR VPWR U$$3691/A sky130_fd_sc_hd__a22o_1
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk _369_/CLK VGND VGND VPWR VPWR _497_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_91_1 dadda_fa_4_91_1/A dadda_fa_4_91_1/B dadda_fa_4_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/B dadda_fa_5_91_1/B sky130_fd_sc_hd__fa_1
XFILLER_181_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_84_0 dadda_fa_4_84_0/A dadda_fa_4_84_0/B dadda_fa_4_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/A dadda_fa_5_84_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_105_3 dadda_fa_3_105_3/A dadda_fa_3_105_3/B dadda_fa_3_105_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_106_1/B dadda_fa_4_105_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_672_ _677_/CLK _672_/D VGND VGND VPWR VPWR _672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$801 U$$938/A1 U$$689/X U$$940/A1 U$$690/X VGND VGND VPWR VPWR U$$802/A sky130_fd_sc_hd__a22o_1
XU$$812 U$$812/A _627_/Q VGND VGND VPWR VPWR U$$812/X sky130_fd_sc_hd__xor2_1
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$823 _628_/Q VGND VGND VPWR VPWR U$$825/B sky130_fd_sc_hd__inv_1
XU$$834 U$$971/A1 U$$928/A2 U$$12/B1 U$$928/B2 VGND VGND VPWR VPWR U$$835/A sky130_fd_sc_hd__a22o_1
XFILLER_21_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$845 U$$845/A U$$923/B VGND VGND VPWR VPWR U$$845/X sky130_fd_sc_hd__xor2_1
XFILLER_90_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$856 U$$34/A1 U$$928/A2 U$$36/A1 U$$928/B2 VGND VGND VPWR VPWR U$$857/A sky130_fd_sc_hd__a22o_1
XU$$867 U$$867/A U$$923/B VGND VGND VPWR VPWR U$$867/X sky130_fd_sc_hd__xor2_1
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1006 U$$1006/A U$$980/B VGND VGND VPWR VPWR U$$1006/X sky130_fd_sc_hd__xor2_1
XU$$1017 U$$58/A1 U$$999/A2 U$$60/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1018/A sky130_fd_sc_hd__a22o_1
XU$$878 U$$878/A1 U$$910/A2 U$$880/A1 U$$910/B2 VGND VGND VPWR VPWR U$$879/A sky130_fd_sc_hd__a22o_1
XU$$889 U$$889/A U$$923/B VGND VGND VPWR VPWR U$$889/X sky130_fd_sc_hd__xor2_1
XU$$1028 U$$1028/A U$$980/B VGND VGND VPWR VPWR U$$1028/X sky130_fd_sc_hd__xor2_1
XU$$1039 U$$902/A1 U$$999/A2 U$$902/B1 U$$987/B2 VGND VGND VPWR VPWR U$$1040/A sky130_fd_sc_hd__a22o_1
XFILLER_189_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _336_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_99_0 dadda_fa_6_99_0/A dadda_fa_6_99_0/B dadda_fa_6_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_100_0/B dadda_fa_7_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_41_4 dadda_fa_2_41_4/A dadda_fa_2_41_4/B dadda_fa_2_41_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_1/CIN dadda_fa_3_41_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_34_3 U$$1538/X U$$1671/X U$$1804/X VGND VGND VPWR VPWR dadda_fa_3_35_1/B
+ dadda_fa_3_34_3/B sky130_fd_sc_hd__fa_1
XFILLER_35_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2230 _567_/Q U$$2196/X U$$3191/A1 U$$2197/X VGND VGND VPWR VPWR U$$2231/A sky130_fd_sc_hd__a22o_1
XU$$2241 U$$2241/A U$$2257/B VGND VGND VPWR VPWR U$$2241/X sky130_fd_sc_hd__xor2_1
XFILLER_35_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2252 U$$4170/A1 U$$2270/A2 U$$3624/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2253/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2263 U$$2263/A U$$2327/B VGND VGND VPWR VPWR U$$2263/X sky130_fd_sc_hd__xor2_1
XFILLER_62_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2274 _589_/Q U$$2326/A2 _590_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2275/A sky130_fd_sc_hd__a22o_1
XU$$1540 U$$1540/A U$$1580/B VGND VGND VPWR VPWR U$$1540/X sky130_fd_sc_hd__xor2_1
XU$$2285 U$$2285/A U$$2289/B VGND VGND VPWR VPWR U$$2285/X sky130_fd_sc_hd__xor2_1
XU$$2296 U$$926/A1 U$$2316/A2 _601_/Q U$$2316/B2 VGND VGND VPWR VPWR U$$2297/A sky130_fd_sc_hd__a22o_1
XU$$1551 U$$4291/A1 U$$1591/A2 U$$868/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1552/A
+ sky130_fd_sc_hd__a22o_1
XU$$1562 U$$1562/A U$$1580/B VGND VGND VPWR VPWR U$$1562/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1573 U$$3489/B1 U$$1605/A2 U$$3217/B1 U$$1605/B2 VGND VGND VPWR VPWR U$$1574/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _331_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1584 U$$1584/A U$$1643/A VGND VGND VPWR VPWR U$$1584/X sky130_fd_sc_hd__xor2_1
XFILLER_176_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1595 U$$771/B1 U$$1511/X U$$90/A1 U$$1512/X VGND VGND VPWR VPWR U$$1596/A sky130_fd_sc_hd__a22o_1
XFILLER_33_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_79_5 U$$3091/X U$$3224/X U$$3357/X VGND VGND VPWR VPWR dadda_fa_2_80_2/A
+ dadda_fa_2_79_5/A sky130_fd_sc_hd__fa_1
XFILLER_98_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$203 final_adder.U$$697/A final_adder.U$$569/B1 final_adder.U$$203/B1
+ VGND VGND VPWR VPWR final_adder.U$$203/X sky130_fd_sc_hd__a21o_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$214 final_adder.U$$709/A final_adder.U$$708/A VGND VGND VPWR VPWR
+ final_adder.U$$298/A sky130_fd_sc_hd__and2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$225 final_adder.U$$719/A final_adder.U$$591/B1 final_adder.U$$225/B1
+ VGND VGND VPWR VPWR final_adder.U$$225/X sky130_fd_sc_hd__a21o_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$236 final_adder.U$$731/A final_adder.U$$730/A VGND VGND VPWR VPWR
+ final_adder.U$$310/B sky130_fd_sc_hd__and2_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater440 U$$1770/A2 VGND VGND VPWR VPWR U$$1726/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$247 final_adder.U$$741/A final_adder.U$$613/B1 final_adder.U$$247/B1
+ VGND VGND VPWR VPWR final_adder.U$$247/X sky130_fd_sc_hd__a21o_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater451 U$$1100/X VGND VGND VPWR VPWR U$$1218/A2 sky130_fd_sc_hd__buf_12
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater462 U$$4115/X VGND VGND VPWR VPWR U$$4198/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$258 final_adder.U$$258/A final_adder.U$$258/B VGND VGND VPWR VPWR
+ final_adder.U$$258/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$269 final_adder.U$$268/A final_adder.U$$153/X final_adder.U$$155/X
+ VGND VGND VPWR VPWR final_adder.U$$269/X sky130_fd_sc_hd__a21o_1
XU$$108 U$$930/A1 U$$4/X _603_/Q U$$5/X VGND VGND VPWR VPWR U$$109/A sky130_fd_sc_hd__a22o_1
Xrepeater473 U$$3430/X VGND VGND VPWR VPWR U$$3545/B2 sky130_fd_sc_hd__buf_12
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$119 U$$119/A U$$3/A VGND VGND VPWR VPWR U$$119/X sky130_fd_sc_hd__xor2_1
Xrepeater484 U$$2745/X VGND VGND VPWR VPWR U$$2870/B2 sky130_fd_sc_hd__buf_12
XFILLER_66_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater495 U$$2189/B2 VGND VGND VPWR VPWR U$$2161/B2 sky130_fd_sc_hd__buf_12
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_110_1 U$$3552/X U$$3685/X U$$3818/X VGND VGND VPWR VPWR dadda_fa_4_111_1/A
+ dadda_fa_4_110_2/A sky130_fd_sc_hd__fa_1
XFILLER_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_0 U$$3937/X U$$4070/X U$$4203/X VGND VGND VPWR VPWR dadda_fa_4_104_0/B
+ dadda_fa_4_103_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_68_5 U$$2271/X U$$2404/X VGND VGND VPWR VPWR dadda_fa_1_69_7/B dadda_fa_2_68_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_49_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput210 c[58] VGND VGND VPWR VPWR input210/X sky130_fd_sc_hd__buf_4
XFILLER_49_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput221 c[68] VGND VGND VPWR VPWR input221/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput232 c[78] VGND VGND VPWR VPWR input232/X sky130_fd_sc_hd__clkbuf_1
Xinput243 c[88] VGND VGND VPWR VPWR input243/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_51_3 dadda_fa_3_51_3/A dadda_fa_3_51_3/B dadda_fa_3_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/B dadda_fa_4_51_2/CIN sky130_fd_sc_hd__fa_1
Xinput254 c[98] VGND VGND VPWR VPWR input254/X sky130_fd_sc_hd__buf_2
Xdadda_fa_0_67_3 U$$1338/X U$$1471/X U$$1604/X VGND VGND VPWR VPWR dadda_fa_1_68_6/B
+ dadda_fa_1_67_8/B sky130_fd_sc_hd__fa_1
XFILLER_64_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_44_2 dadda_fa_3_44_2/A dadda_fa_3_44_2/B dadda_fa_3_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/A dadda_fa_4_44_2/B sky130_fd_sc_hd__fa_1
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_37_1 dadda_fa_3_37_1/A dadda_fa_3_37_1/B dadda_fa_3_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/CIN dadda_fa_4_37_2/A sky130_fd_sc_hd__fa_2
XU$$620 U$$70/B1 U$$626/A2 U$$759/A1 U$$553/X VGND VGND VPWR VPWR U$$621/A sky130_fd_sc_hd__a22o_1
XFILLER_29_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$631 U$$631/A U$$661/B VGND VGND VPWR VPWR U$$631/X sky130_fd_sc_hd__xor2_1
X_655_ _667_/CLK _655_/D VGND VGND VPWR VPWR _655_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$642 U$$92/B1 U$$682/A2 U$$96/A1 U$$553/X VGND VGND VPWR VPWR U$$643/A sky130_fd_sc_hd__a22o_1
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_14_0 dadda_fa_6_14_0/A dadda_fa_6_14_0/B dadda_fa_6_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_15_0/B dadda_fa_7_14_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$653 U$$653/A U$$661/B VGND VGND VPWR VPWR U$$653/X sky130_fd_sc_hd__xor2_1
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$664 U$$938/A1 U$$552/X U$$940/A1 U$$553/X VGND VGND VPWR VPWR U$$665/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$675 U$$675/A _625_/Q VGND VGND VPWR VPWR U$$675/X sky130_fd_sc_hd__xor2_1
XU$$686 _626_/Q VGND VGND VPWR VPWR U$$688/B sky130_fd_sc_hd__inv_1
X_586_ _679_/CLK _586_/D VGND VGND VPWR VPWR _586_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_90_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$697 U$$971/A1 U$$817/A2 U$$12/B1 U$$785/B2 VGND VGND VPWR VPWR U$$698/A sky130_fd_sc_hd__a22o_1
XFILLER_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_96_5 U$$4455/X input252/X dadda_fa_2_96_5/CIN VGND VGND VPWR VPWR dadda_fa_3_97_2/A
+ dadda_fa_4_96_0/A sky130_fd_sc_hd__fa_2
XFILLER_181_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_89_4 dadda_fa_2_89_4/A dadda_fa_2_89_4/B dadda_fa_2_89_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_1/CIN dadda_fa_3_89_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_193_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_clk _431_/CLK VGND VGND VPWR VPWR _327_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_32_0 U$$71/X U$$204/X U$$337/X VGND VGND VPWR VPWR dadda_fa_3_33_0/B dadda_fa_3_32_2/B
+ sky130_fd_sc_hd__fa_2
XFILLER_82_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2060 U$$2058/B U$$2055/A _646_/Q U$$2055/Y VGND VGND VPWR VPWR U$$2060/X sky130_fd_sc_hd__a22o_4
XU$$2071 U$$14/B1 U$$2117/A2 U$$4265/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2072/A sky130_fd_sc_hd__a22o_1
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2082 U$$2082/A U$$2118/B VGND VGND VPWR VPWR U$$2082/X sky130_fd_sc_hd__xor2_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2093 U$$4285/A1 U$$2117/A2 U$$3191/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2094/A
+ sky130_fd_sc_hd__a22o_1
XU$$1370 _635_/Q VGND VGND VPWR VPWR U$$1370/Y sky130_fd_sc_hd__inv_1
XU$$1381 U$$1381/A U$$1479/B VGND VGND VPWR VPWR U$$1381/X sky130_fd_sc_hd__xor2_1
XFILLER_149_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1392 U$$979/B1 U$$1472/A2 U$$983/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1393/A sky130_fd_sc_hd__a22o_1
XFILLER_176_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_119_0 input150/X dadda_fa_5_119_0/B dadda_fa_5_119_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_6_120_0/A dadda_fa_6_119_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_84_3 U$$2569/X U$$2702/X U$$2835/X VGND VGND VPWR VPWR dadda_fa_2_85_3/A
+ dadda_fa_2_84_5/A sky130_fd_sc_hd__fa_1
XFILLER_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_61_2 dadda_fa_4_61_2/A dadda_fa_4_61_2/B dadda_fa_4_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/CIN dadda_fa_5_61_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_77_2 U$$2156/X U$$2289/X U$$2422/X VGND VGND VPWR VPWR dadda_fa_2_78_1/A
+ dadda_fa_2_77_4/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_54_1 dadda_fa_4_54_1/A dadda_fa_4_54_1/B dadda_fa_4_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/B dadda_fa_5_54_1/B sky130_fd_sc_hd__fa_1
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_31_0 dadda_fa_7_31_0/A dadda_fa_7_31_0/B dadda_fa_7_31_0/CIN VGND VGND
+ VPWR VPWR _456_/D _327_/D sky130_fd_sc_hd__fa_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_47_0 dadda_fa_4_47_0/A dadda_fa_4_47_0/B dadda_fa_4_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/A dadda_fa_5_47_1/A sky130_fd_sc_hd__fa_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _463_/CLK _440_/D VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _500_/CLK _371_/D VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_99_3 dadda_fa_3_99_3/A dadda_fa_3_99_3/B dadda_fa_3_99_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/B dadda_fa_4_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_72_1 U$$949/X U$$1082/X U$$1215/X VGND VGND VPWR VPWR dadda_fa_1_73_7/B
+ dadda_fa_1_72_8/B sky130_fd_sc_hd__fa_1
XFILLER_89_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_65_0 U$$89/B U$$270/X U$$403/X VGND VGND VPWR VPWR dadda_fa_1_66_5/B dadda_fa_1_65_7/B
+ sky130_fd_sc_hd__fa_1
XFILLER_37_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$450 U$$450/A U$$530/B VGND VGND VPWR VPWR U$$450/X sky130_fd_sc_hd__xor2_1
XFILLER_189_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_638_ _642_/CLK _638_/D VGND VGND VPWR VPWR _638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$461 U$$735/A1 U$$545/A2 U$$52/A1 U$$416/X VGND VGND VPWR VPWR U$$462/A sky130_fd_sc_hd__a22o_1
XU$$472 U$$472/A U$$547/A VGND VGND VPWR VPWR U$$472/X sky130_fd_sc_hd__xor2_1
XFILLER_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$483 U$$72/A1 U$$491/A2 U$$74/A1 U$$416/X VGND VGND VPWR VPWR U$$484/A sky130_fd_sc_hd__a22o_1
XU$$494 U$$494/A _623_/Q VGND VGND VPWR VPWR U$$494/X sky130_fd_sc_hd__xor2_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_569_ _576_/CLK _569_/D VGND VGND VPWR VPWR _569_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_94_2 U$$3520/X U$$3653/X U$$3786/X VGND VGND VPWR VPWR dadda_fa_3_95_1/A
+ dadda_fa_3_94_3/A sky130_fd_sc_hd__fa_2
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_71_1 dadda_fa_5_71_1/A dadda_fa_5_71_1/B dadda_fa_5_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/B dadda_fa_7_71_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_87_1 U$$4038/X U$$4171/X U$$4304/X VGND VGND VPWR VPWR dadda_fa_3_88_0/CIN
+ dadda_fa_3_87_2/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_5_64_0 dadda_fa_5_64_0/A dadda_fa_5_64_0/B dadda_fa_5_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/A dadda_fa_6_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_63_8 dadda_fa_1_63_8/A dadda_fa_1_63_8/B dadda_fa_1_63_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_3/A dadda_fa_3_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_56_7 U$$3893/B input208/X dadda_fa_1_56_7/CIN VGND VGND VPWR VPWR dadda_fa_2_57_2/CIN
+ dadda_fa_2_56_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_49_6 U$$2499/X U$$2632/X U$$2765/X VGND VGND VPWR VPWR dadda_fa_2_50_2/CIN
+ dadda_fa_2_49_5/CIN sky130_fd_sc_hd__fa_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_90_3 U$$2980/X U$$3113/X VGND VGND VPWR VPWR dadda_fa_2_91_5/A dadda_fa_3_90_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_79_0 dadda_fa_7_79_0/A dadda_fa_7_79_0/B dadda_fa_7_79_0/CIN VGND VGND
+ VPWR VPWR _504_/D _375_/D sky130_fd_sc_hd__fa_1
XFILLER_108_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_82_0 _686__906/HI U$$1368/X U$$1501/X VGND VGND VPWR VPWR dadda_fa_2_83_1/B
+ dadda_fa_2_82_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_132_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4209 U$$4209/A _677_/Q VGND VGND VPWR VPWR U$$4209/X sky130_fd_sc_hd__xor2_1
XFILLER_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3508 U$$3508/A U$$3536/B VGND VGND VPWR VPWR U$$3508/X sky130_fd_sc_hd__xor2_1
XFILLER_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3519 U$$94/A1 U$$3429/X U$$94/B1 U$$3430/X VGND VGND VPWR VPWR U$$3520/A sky130_fd_sc_hd__a22o_1
XFILLER_18_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2807 U$$2807/A U$$2839/B VGND VGND VPWR VPWR U$$2807/X sky130_fd_sc_hd__xor2_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2818 U$$76/B1 U$$2868/A2 U$$902/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2819/A sky130_fd_sc_hd__a22o_1
XU$$2829 U$$2829/A U$$2871/B VGND VGND VPWR VPWR U$$2829/X sky130_fd_sc_hd__xor2_1
XFILLER_65_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _551_/CLK _423_/D VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_354_ _490_/CLK _354_/D VGND VGND VPWR VPWR _354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_285_ _612_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_81_0 dadda_fa_6_81_0/A dadda_fa_6_81_0/B dadda_fa_6_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_82_0/B dadda_fa_7_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_97_0 dadda_fa_3_97_0/A dadda_fa_3_97_0/B dadda_fa_3_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/B dadda_fa_4_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_182_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_59_5 dadda_fa_2_59_5/A dadda_fa_2_59_5/B dadda_fa_2_59_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_2/A dadda_fa_4_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput7 a[15] VGND VGND VPWR VPWR _631_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_92_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$280 U$$280/A1 U$$278/X U$$8/A1 U$$279/X VGND VGND VPWR VPWR U$$281/A sky130_fd_sc_hd__a22o_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$291 U$$291/A U$$391/B VGND VGND VPWR VPWR U$$291/X sky130_fd_sc_hd__xor2_1
XFILLER_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$5 _429_/Q _301_/Q VGND VGND VPWR VPWR final_adder.U$$5/COUT final_adder.U$$627/A
+ sky130_fd_sc_hd__ha_2
Xoutput300 _191_/Q VGND VGND VPWR VPWR o[23] sky130_fd_sc_hd__buf_2
Xoutput311 _201_/Q VGND VGND VPWR VPWR o[33] sky130_fd_sc_hd__buf_2
XFILLER_160_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput322 _211_/Q VGND VGND VPWR VPWR o[43] sky130_fd_sc_hd__buf_2
XFILLER_161_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput333 _221_/Q VGND VGND VPWR VPWR o[53] sky130_fd_sc_hd__buf_2
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput344 _231_/Q VGND VGND VPWR VPWR o[63] sky130_fd_sc_hd__buf_2
Xoutput355 _241_/Q VGND VGND VPWR VPWR o[73] sky130_fd_sc_hd__buf_2
XFILLER_142_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput366 _251_/Q VGND VGND VPWR VPWR o[83] sky130_fd_sc_hd__buf_2
Xoutput377 _261_/Q VGND VGND VPWR VPWR o[93] sky130_fd_sc_hd__buf_2
XFILLER_160_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_61_5 U$$3986/X U$$4119/X input214/X VGND VGND VPWR VPWR dadda_fa_2_62_2/A
+ dadda_fa_2_61_5/A sky130_fd_sc_hd__fa_2
XFILLER_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_54_4 U$$2376/X U$$2509/X U$$2642/X VGND VGND VPWR VPWR dadda_fa_2_55_1/CIN
+ dadda_fa_2_54_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_47_3 U$$1298/X U$$1431/X U$$1564/X VGND VGND VPWR VPWR dadda_fa_2_48_2/B
+ dadda_fa_2_47_5/A sky130_fd_sc_hd__fa_1
XFILLER_56_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_24_2 dadda_fa_4_24_2/A dadda_fa_4_24_2/B dadda_fa_4_24_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/CIN dadda_fa_5_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_1 U$$1105/X input165/X dadda_fa_4_17_1/CIN VGND VGND VPWR VPWR dadda_fa_5_18_0/B
+ dadda_fa_5_17_1/B sky130_fd_sc_hd__fa_1
XFILLER_169_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4006 U$$4006/A U$$4058/B VGND VGND VPWR VPWR U$$4006/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_20_3 U$$1244/X U$$1377/X VGND VGND VPWR VPWR dadda_fa_4_21_1/B dadda_ha_3_20_3/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4017 U$$4289/B1 U$$3977/X U$$4291/B1 U$$3978/X VGND VGND VPWR VPWR U$$4018/A sky130_fd_sc_hd__a22o_1
XFILLER_120_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4028 U$$4028/A U$$4044/B VGND VGND VPWR VPWR U$$4028/X sky130_fd_sc_hd__xor2_1
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4039 _581_/Q U$$4045/A2 U$$4178/A1 U$$3978/X VGND VGND VPWR VPWR U$$4040/A sky130_fd_sc_hd__a22o_1
XU$$3305 U$$3305/A U$$3397/B VGND VGND VPWR VPWR U$$3305/X sky130_fd_sc_hd__xor2_1
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3316 _562_/Q U$$3396/A2 _563_/Q U$$3396/B2 VGND VGND VPWR VPWR U$$3317/A sky130_fd_sc_hd__a22o_1
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3327 U$$3327/A U$$3413/B VGND VGND VPWR VPWR U$$3327/X sky130_fd_sc_hd__xor2_1
XFILLER_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3338 _573_/Q U$$3396/A2 U$$50/B1 U$$3396/B2 VGND VGND VPWR VPWR U$$3339/A sky130_fd_sc_hd__a22o_1
XU$$2604 _654_/Q VGND VGND VPWR VPWR U$$2606/B sky130_fd_sc_hd__inv_1
XU$$3349 U$$3349/A U$$3397/B VGND VGND VPWR VPWR U$$3349/X sky130_fd_sc_hd__xor2_1
XU$$2615 U$$12/A1 U$$2729/A2 _555_/Q U$$2729/B2 VGND VGND VPWR VPWR U$$2616/A sky130_fd_sc_hd__a22o_1
XU$$2626 U$$2626/A U$$2694/B VGND VGND VPWR VPWR U$$2626/X sky130_fd_sc_hd__xor2_1
XFILLER_62_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2637 _565_/Q U$$2667/A2 U$$4283/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2638/A sky130_fd_sc_hd__a22o_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2648 U$$2648/A U$$2698/B VGND VGND VPWR VPWR U$$2648/X sky130_fd_sc_hd__xor2_1
XU$$1903 _609_/Q U$$1903/A2 _610_/Q U$$1903/B2 VGND VGND VPWR VPWR U$$1904/A sky130_fd_sc_hd__a22o_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1914 U$$1914/A _643_/Q VGND VGND VPWR VPWR U$$1914/X sky130_fd_sc_hd__xor2_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2659 U$$878/A1 U$$2667/A2 U$$880/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2660/A sky130_fd_sc_hd__a22o_1
XU$$1925 U$$1925/A U$$2021/B VGND VGND VPWR VPWR U$$1925/X sky130_fd_sc_hd__xor2_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1936 U$$4265/A1 U$$2036/A2 U$$979/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$1937/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1947 U$$1947/A U$$2021/B VGND VGND VPWR VPWR U$$1947/X sky130_fd_sc_hd__xor2_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1958 U$$3191/A1 U$$2048/A2 U$$3876/B1 U$$2048/B2 VGND VGND VPWR VPWR U$$1959/A
+ sky130_fd_sc_hd__a22o_1
X_406_ _543_/CLK _406_/D VGND VGND VPWR VPWR _406_/Q sky130_fd_sc_hd__dfxtp_1
XU$$1969 U$$1969/A U$$2021/B VGND VGND VPWR VPWR U$$1969/X sky130_fd_sc_hd__xor2_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_337_ _467_/CLK _337_/D VGND VGND VPWR VPWR _337_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ _280_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_199_ _329_/CLK _199_/D VGND VGND VPWR VPWR _199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_4 dadda_fa_2_71_4/A dadda_fa_2_71_4/B dadda_fa_2_71_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/CIN dadda_fa_3_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_64_3 dadda_fa_2_64_3/A dadda_fa_2_64_3/B dadda_fa_2_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/B dadda_fa_3_64_3/B sky130_fd_sc_hd__fa_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_1_1_1_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_57_2 dadda_fa_2_57_2/A dadda_fa_2_57_2/B dadda_fa_2_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/A dadda_fa_3_57_3/A sky130_fd_sc_hd__fa_2
XU$$10 U$$8/B1 U$$4/X U$$12/A1 U$$5/X VGND VGND VPWR VPWR U$$11/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_34_1 dadda_fa_5_34_1/A dadda_fa_5_34_1/B dadda_fa_5_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/B dadda_fa_7_34_0/A sky130_fd_sc_hd__fa_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$21 U$$21/A U$$9/B VGND VGND VPWR VPWR U$$21/X sky130_fd_sc_hd__xor2_1
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$32 U$$32/A1 U$$4/X U$$34/A1 U$$5/X VGND VGND VPWR VPWR U$$33/A sky130_fd_sc_hd__a22o_1
XU$$43 U$$43/A U$$3/A VGND VGND VPWR VPWR U$$43/X sky130_fd_sc_hd__xor2_1
XFILLER_53_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$54 U$$54/A1 U$$4/X U$$56/A1 U$$5/X VGND VGND VPWR VPWR U$$55/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_27_0 dadda_fa_5_27_0/A dadda_fa_5_27_0/B dadda_fa_5_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/A dadda_fa_6_27_0/CIN sky130_fd_sc_hd__fa_1
XU$$3850 U$$14/A1 U$$3840/X _556_/Q U$$3841/X VGND VGND VPWR VPWR U$$3851/A sky130_fd_sc_hd__a22o_1
XU$$65 U$$65/A U$$89/B VGND VGND VPWR VPWR U$$65/X sky130_fd_sc_hd__xor2_1
XU$$3861 U$$3861/A U$$3893/B VGND VGND VPWR VPWR U$$3861/X sky130_fd_sc_hd__xor2_1
XU$$76 U$$76/A1 U$$4/X U$$76/B1 U$$5/X VGND VGND VPWR VPWR U$$77/A sky130_fd_sc_hd__a22o_1
XU$$3872 U$$4283/A1 U$$3840/X U$$4285/A1 U$$3841/X VGND VGND VPWR VPWR U$$3873/A sky130_fd_sc_hd__a22o_1
XU$$87 U$$87/A U$$3/A VGND VGND VPWR VPWR U$$87/X sky130_fd_sc_hd__xor2_1
XFILLER_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3883 U$$3883/A U$$3969/B VGND VGND VPWR VPWR U$$3883/X sky130_fd_sc_hd__xor2_1
XU$$98 U$$98/A1 U$$4/X U$$98/B1 U$$5/X VGND VGND VPWR VPWR U$$99/A sky130_fd_sc_hd__a22o_1
XU$$3894 _577_/Q U$$3912/A2 U$$4170/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3895/A sky130_fd_sc_hd__a22o_1
XFILLER_75_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_101_0 dadda_fa_5_101_0/A dadda_fa_5_101_0/B dadda_fa_5_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/A dadda_fa_6_101_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_830__882 VGND VGND VPWR VPWR _830__882/HI U$$4505/B sky130_fd_sc_hd__conb_1
XFILLER_133_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_52_1 U$$776/X U$$909/X U$$1042/X VGND VGND VPWR VPWR dadda_fa_2_53_0/CIN
+ dadda_fa_2_52_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_45_0 U$$97/X U$$230/X U$$363/X VGND VGND VPWR VPWR dadda_fa_2_46_2/A dadda_fa_2_45_4/B
+ sky130_fd_sc_hd__fa_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_81_3 dadda_fa_3_81_3/A dadda_fa_3_81_3/B dadda_fa_3_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/B dadda_fa_4_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_74_2 dadda_fa_3_74_2/A dadda_fa_3_74_2/B dadda_fa_3_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/A dadda_fa_4_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_67_1 dadda_fa_3_67_1/A dadda_fa_3_67_1/B dadda_fa_3_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/CIN dadda_fa_4_67_2/A sky130_fd_sc_hd__fa_1
XFILLER_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_44_0 dadda_fa_6_44_0/A dadda_fa_6_44_0/B dadda_fa_6_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_45_0/B dadda_fa_7_44_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3102 U$$771/B1 U$$3018/X U$$912/A1 U$$3019/X VGND VGND VPWR VPWR U$$3103/A sky130_fd_sc_hd__a22o_1
XU$$3113 U$$3113/A U$$3137/B VGND VGND VPWR VPWR U$$3113/X sky130_fd_sc_hd__xor2_1
XU$$3124 _603_/Q U$$3018/X _604_/Q U$$3019/X VGND VGND VPWR VPWR U$$3125/A sky130_fd_sc_hd__a22o_1
XFILLER_19_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3135 U$$3135/A U$$3137/B VGND VGND VPWR VPWR U$$3135/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2401 U$$70/B1 U$$2333/X U$$759/A1 U$$2334/X VGND VGND VPWR VPWR U$$2402/A sky130_fd_sc_hd__a22o_1
XU$$3146 U$$4379/A1 U$$3146/A2 U$$956/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3147/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2412 U$$2412/A U$$2436/B VGND VGND VPWR VPWR U$$2412/X sky130_fd_sc_hd__xor2_1
XU$$3157 U$$3157/A1 U$$3241/A2 U$$4255/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3158/A
+ sky130_fd_sc_hd__a22o_1
XU$$2423 _595_/Q U$$2463/A2 _596_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2424/A sky130_fd_sc_hd__a22o_1
XU$$3168 U$$3168/A U$$3244/B VGND VGND VPWR VPWR U$$3168/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_2 dadda_fa_4_103_2/A dadda_fa_4_103_2/B dadda_fa_4_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/CIN dadda_fa_5_103_1/CIN sky130_fd_sc_hd__fa_1
XU$$2434 U$$2434/A U$$2436/B VGND VGND VPWR VPWR U$$2434/X sky130_fd_sc_hd__xor2_1
XFILLER_35_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3179 U$$28/A1 U$$3241/A2 U$$30/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3180/A sky130_fd_sc_hd__a22o_1
XU$$2445 _606_/Q U$$2463/A2 U$$940/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2446/A sky130_fd_sc_hd__a22o_1
XU$$1700 U$$878/A1 U$$1726/A2 U$$880/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1701/A sky130_fd_sc_hd__a22o_1
XU$$1711 U$$1711/A U$$1739/B VGND VGND VPWR VPWR U$$1711/X sky130_fd_sc_hd__xor2_1
XU$$2456 U$$2456/A U$$2464/B VGND VGND VPWR VPWR U$$2456/X sky130_fd_sc_hd__xor2_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2467 _652_/Q VGND VGND VPWR VPWR U$$2469/B sky130_fd_sc_hd__inv_1
XU$$1722 U$$76/B1 U$$1770/A2 U$$902/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1723/A sky130_fd_sc_hd__a22o_1
XFILLER_185_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1733 U$$1733/A U$$1781/A VGND VGND VPWR VPWR U$$1733/X sky130_fd_sc_hd__xor2_1
XFILLER_15_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2478 U$$971/A1 U$$2574/A2 U$$12/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2479/A sky130_fd_sc_hd__a22o_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2489 U$$2489/A U$$2533/B VGND VGND VPWR VPWR U$$2489/X sky130_fd_sc_hd__xor2_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1744 _598_/Q U$$1770/A2 _599_/Q U$$1770/B2 VGND VGND VPWR VPWR U$$1745/A sky130_fd_sc_hd__a22o_1
XU$$1755 U$$1755/A U$$1781/A VGND VGND VPWR VPWR U$$1755/X sky130_fd_sc_hd__xor2_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1766 U$$944/A1 U$$1648/X U$$946/A1 U$$1649/X VGND VGND VPWR VPWR U$$1767/A sky130_fd_sc_hd__a22o_1
XFILLER_187_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1777 U$$1777/A _641_/Q VGND VGND VPWR VPWR U$$1777/X sky130_fd_sc_hd__xor2_1
XU$$1788 U$$1788/A U$$1918/A VGND VGND VPWR VPWR U$$1788/X sky130_fd_sc_hd__xor2_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1799 U$$18/A1 U$$1867/A2 U$$20/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1800/A sky130_fd_sc_hd__a22o_1
XFILLER_188_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_773__825 VGND VGND VPWR VPWR _773__825/HI U$$4391/B sky130_fd_sc_hd__conb_1
Xdadda_fa_7_117_0 dadda_fa_7_117_0/A dadda_fa_7_117_0/B dadda_fa_7_117_0/CIN VGND
+ VGND VPWR VPWR _542_/D _413_/D sky130_fd_sc_hd__fa_2
Xinput10 a[18] VGND VGND VPWR VPWR _634_/D sky130_fd_sc_hd__buf_2
Xinput21 a[28] VGND VGND VPWR VPWR _644_/D sky130_fd_sc_hd__buf_2
Xinput32 a[38] VGND VGND VPWR VPWR _654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput43 a[48] VGND VGND VPWR VPWR _664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput54 a[58] VGND VGND VPWR VPWR _674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput65 b[0] VGND VGND VPWR VPWR _552_/D sky130_fd_sc_hd__buf_2
XFILLER_157_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput76 b[1] VGND VGND VPWR VPWR _553_/D sky130_fd_sc_hd__buf_2
X_814__866 VGND VGND VPWR VPWR _814__866/HI U$$4473/B sky130_fd_sc_hd__conb_1
Xinput87 b[2] VGND VGND VPWR VPWR _554_/D sky130_fd_sc_hd__buf_2
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput98 b[3] VGND VGND VPWR VPWR _555_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_115_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater600 _625_/Q VGND VGND VPWR VPWR U$$623/B sky130_fd_sc_hd__buf_12
XFILLER_85_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_62_0 dadda_fa_2_62_0/A dadda_fa_2_62_0/B dadda_fa_2_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/B dadda_fa_3_62_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$407 final_adder.U$$324/B final_adder.U$$638/B final_adder.U$$265/X
+ VGND VGND VPWR VPWR final_adder.U$$642/B sky130_fd_sc_hd__a21o_1
Xrepeater611 _617_/Q VGND VGND VPWR VPWR U$$89/B sky130_fd_sc_hd__buf_12
XFILLER_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater622 U$$4508/A1 VGND VGND VPWR VPWR U$$946/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$429 final_adder.U$$346/B final_adder.U$$726/B final_adder.U$$309/X
+ VGND VGND VPWR VPWR final_adder.U$$730/B sky130_fd_sc_hd__a21o_1
Xrepeater633 _605_/Q VGND VGND VPWR VPWR U$$799/A1 sky130_fd_sc_hd__buf_12
XFILLER_85_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater644 _600_/Q VGND VGND VPWR VPWR U$$787/B1 sky130_fd_sc_hd__buf_12
Xrepeater655 _595_/Q VGND VGND VPWR VPWR U$$94/A1 sky130_fd_sc_hd__buf_12
Xrepeater666 _591_/Q VGND VGND VPWR VPWR U$$908/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater677 U$$76/A1 VGND VGND VPWR VPWR U$$2953/A1 sky130_fd_sc_hd__buf_12
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater688 _583_/Q VGND VGND VPWR VPWR U$$70/A1 sky130_fd_sc_hd__buf_12
XU$$4370 U$$4370/A U$$4384/A VGND VGND VPWR VPWR U$$4370/X sky130_fd_sc_hd__xor2_1
Xrepeater699 _578_/Q VGND VGND VPWR VPWR U$$60/A1 sky130_fd_sc_hd__buf_12
XU$$4381 U$$819/A1 U$$4381/A2 U$$4381/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4382/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4392 _552_/Q U$$4388/X _553_/Q U$$4389/X VGND VGND VPWR VPWR U$$4393/A sky130_fd_sc_hd__a22o_1
XFILLER_26_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3680 U$$4502/A1 U$$3566/X U$$4504/A1 U$$3567/X VGND VGND VPWR VPWR U$$3681/A sky130_fd_sc_hd__a22o_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3691 U$$3691/A U$$3698/A VGND VGND VPWR VPWR U$$3691/X sky130_fd_sc_hd__xor2_1
XU$$2990 U$$2990/A U$$3004/B VGND VGND VPWR VPWR U$$2990/X sky130_fd_sc_hd__xor2_1
XFILLER_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_91_2 dadda_fa_4_91_2/A dadda_fa_4_91_2/B dadda_fa_4_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/CIN dadda_fa_5_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_10_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_84_1 dadda_fa_4_84_1/A dadda_fa_4_84_1/B dadda_fa_4_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/B dadda_fa_5_84_1/B sky130_fd_sc_hd__fa_1
XFILLER_161_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_61_0 dadda_fa_7_61_0/A dadda_fa_7_61_0/B dadda_fa_7_61_0/CIN VGND VGND
+ VPWR VPWR _486_/D _357_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_77_0 dadda_fa_4_77_0/A dadda_fa_4_77_0/B dadda_fa_4_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/A dadda_fa_5_77_1/A sky130_fd_sc_hd__fa_1
XFILLER_122_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_671_ _679_/CLK _671_/D VGND VGND VPWR VPWR _671_/Q sky130_fd_sc_hd__dfxtp_4
XU$$802 U$$802/A U$$822/A VGND VGND VPWR VPWR U$$802/X sky130_fd_sc_hd__xor2_1
XFILLER_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$813 U$$950/A1 U$$817/A2 U$$952/A1 U$$817/B2 VGND VGND VPWR VPWR U$$814/A sky130_fd_sc_hd__a22o_1
XU$$824 U$$959/A VGND VGND VPWR VPWR U$$824/Y sky130_fd_sc_hd__inv_1
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$835 U$$835/A U$$959/A VGND VGND VPWR VPWR U$$835/X sky130_fd_sc_hd__xor2_1
XFILLER_17_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$846 U$$983/A1 U$$910/A2 U$$26/A1 U$$910/B2 VGND VGND VPWR VPWR U$$847/A sky130_fd_sc_hd__a22o_1
XU$$857 U$$857/A U$$923/B VGND VGND VPWR VPWR U$$857/X sky130_fd_sc_hd__xor2_1
XFILLER_71_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1007 U$$48/A1 U$$999/A2 U$$50/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1008/A sky130_fd_sc_hd__a22o_1
XU$$868 U$$868/A1 U$$910/A2 U$$48/A1 U$$910/B2 VGND VGND VPWR VPWR U$$869/A sky130_fd_sc_hd__a22o_1
XFILLER_113_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1018 U$$1018/A U$$992/B VGND VGND VPWR VPWR U$$1018/X sky130_fd_sc_hd__xor2_1
XU$$879 U$$879/A U$$903/B VGND VGND VPWR VPWR U$$879/X sky130_fd_sc_hd__xor2_1
XU$$1029 U$$68/B1 U$$999/A2 U$$72/A1 U$$987/B2 VGND VGND VPWR VPWR U$$1030/A sky130_fd_sc_hd__a22o_1
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_757__809 VGND VGND VPWR VPWR _757__809/HI U$$3970/B1 sky130_fd_sc_hd__conb_1
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_41_5 dadda_fa_2_41_5/A dadda_fa_2_41_5/B dadda_fa_2_41_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_2/A dadda_fa_4_41_0/A sky130_fd_sc_hd__fa_2
XFILLER_93_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_34_4 U$$1937/X U$$2070/X U$$2203/X VGND VGND VPWR VPWR dadda_fa_3_35_1/CIN
+ dadda_fa_3_34_3/CIN sky130_fd_sc_hd__fa_2
XU$$2220 U$$987/A1 U$$2270/A2 U$$30/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2221/A sky130_fd_sc_hd__a22o_1
XFILLER_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2231 U$$2231/A U$$2289/B VGND VGND VPWR VPWR U$$2231/X sky130_fd_sc_hd__xor2_1
XU$$2242 U$$50/A1 U$$2270/A2 U$$2790/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2243/A sky130_fd_sc_hd__a22o_1
XU$$2253 U$$2253/A U$$2289/B VGND VGND VPWR VPWR U$$2253/X sky130_fd_sc_hd__xor2_1
XU$$2264 U$$70/B1 U$$2196/X U$$759/A1 U$$2197/X VGND VGND VPWR VPWR U$$2265/A sky130_fd_sc_hd__a22o_1
XU$$1530 U$$1530/A U$$1614/B VGND VGND VPWR VPWR U$$1530/X sky130_fd_sc_hd__xor2_1
XFILLER_62_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2275 U$$2275/A U$$2289/B VGND VGND VPWR VPWR U$$2275/X sky130_fd_sc_hd__xor2_1
XU$$1541 U$$3457/B1 U$$1591/A2 U$$4283/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1542/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2286 U$$92/B1 U$$2316/A2 U$$96/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2287/A sky130_fd_sc_hd__a22o_1
XFILLER_22_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2297 U$$2297/A U$$2327/B VGND VGND VPWR VPWR U$$2297/X sky130_fd_sc_hd__xor2_1
XU$$1552 U$$1552/A U$$1580/B VGND VGND VPWR VPWR U$$1552/X sky130_fd_sc_hd__xor2_1
XU$$1563 U$$878/A1 U$$1591/A2 U$$58/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1564/A sky130_fd_sc_hd__a22o_1
XU$$1574 U$$1574/A U$$1580/B VGND VGND VPWR VPWR U$$1574/X sky130_fd_sc_hd__xor2_1
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1585 _587_/Q U$$1605/A2 U$$902/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1586/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1596 U$$1596/A _639_/Q VGND VGND VPWR VPWR U$$1596/X sky130_fd_sc_hd__xor2_1
XFILLER_175_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_94_0 dadda_fa_5_94_0/A dadda_fa_5_94_0/B dadda_fa_5_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/A dadda_fa_6_94_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_79_6 U$$3490/X U$$3623/X U$$3756/X VGND VGND VPWR VPWR dadda_fa_2_80_2/B
+ dadda_fa_2_79_5/B sky130_fd_sc_hd__fa_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$204 final_adder.U$$699/A final_adder.U$$698/A VGND VGND VPWR VPWR
+ final_adder.U$$294/B sky130_fd_sc_hd__and2_1
XFILLER_57_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$215 final_adder.U$$709/A final_adder.U$$581/B1 final_adder.U$$215/B1
+ VGND VGND VPWR VPWR final_adder.U$$215/X sky130_fd_sc_hd__a21o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$226 final_adder.U$$721/A final_adder.U$$720/A VGND VGND VPWR VPWR
+ final_adder.U$$304/A sky130_fd_sc_hd__and2_1
Xrepeater430 U$$2196/X VGND VGND VPWR VPWR U$$2316/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$237 final_adder.U$$731/A final_adder.U$$603/B1 final_adder.U$$237/B1
+ VGND VGND VPWR VPWR final_adder.U$$237/X sky130_fd_sc_hd__a21o_1
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater441 U$$1770/A2 VGND VGND VPWR VPWR U$$1734/A2 sky130_fd_sc_hd__buf_12
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$248 final_adder.U$$743/A final_adder.U$$742/A VGND VGND VPWR VPWR
+ final_adder.U$$316/B sky130_fd_sc_hd__and2_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater452 U$$1073/B2 VGND VGND VPWR VPWR U$$987/B2 sky130_fd_sc_hd__buf_12
Xrepeater463 U$$4063/B2 VGND VGND VPWR VPWR U$$4107/B2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$259 final_adder.U$$258/A final_adder.U$$133/X final_adder.U$$135/X
+ VGND VGND VPWR VPWR final_adder.U$$259/X sky130_fd_sc_hd__a21o_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$109 U$$109/A U$$3/A VGND VGND VPWR VPWR U$$109/X sky130_fd_sc_hd__xor2_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater474 U$$3293/X VGND VGND VPWR VPWR U$$3396/B2 sky130_fd_sc_hd__buf_12
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater485 U$$2729/B2 VGND VGND VPWR VPWR U$$2667/B2 sky130_fd_sc_hd__buf_12
Xrepeater496 U$$2060/X VGND VGND VPWR VPWR U$$2189/B2 sky130_fd_sc_hd__buf_12
XFILLER_72_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_110_2 U$$3951/X U$$4084/X U$$4217/X VGND VGND VPWR VPWR dadda_fa_4_111_1/B
+ dadda_fa_4_110_2/B sky130_fd_sc_hd__fa_1
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_1 U$$4336/X U$$4469/X input133/X VGND VGND VPWR VPWR dadda_fa_4_104_0/CIN
+ dadda_fa_4_103_2/A sky130_fd_sc_hd__fa_2
XFILLER_49_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput200 c[49] VGND VGND VPWR VPWR input200/X sky130_fd_sc_hd__buf_2
Xinput211 c[59] VGND VGND VPWR VPWR input211/X sky130_fd_sc_hd__buf_2
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_124_0 dadda_fa_6_124_0/A dadda_fa_6_124_0/B dadda_fa_6_124_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_125_0/B dadda_fa_7_124_0/CIN sky130_fd_sc_hd__fa_1
Xinput222 c[69] VGND VGND VPWR VPWR input222/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput233 c[79] VGND VGND VPWR VPWR input233/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput244 c[89] VGND VGND VPWR VPWR input244/X sky130_fd_sc_hd__buf_2
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput255 c[99] VGND VGND VPWR VPWR input255/X sky130_fd_sc_hd__buf_2
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_67_4 U$$1737/X U$$1870/X U$$2003/X VGND VGND VPWR VPWR dadda_fa_1_68_6/CIN
+ dadda_fa_1_67_8/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_44_3 dadda_fa_3_44_3/A dadda_fa_3_44_3/B dadda_fa_3_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/B dadda_fa_4_44_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_57_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_654_ _656_/CLK _654_/D VGND VGND VPWR VPWR _654_/Q sky130_fd_sc_hd__dfxtp_1
XU$$610 U$$62/A1 U$$682/A2 U$$64/A1 U$$553/X VGND VGND VPWR VPWR U$$611/A sky130_fd_sc_hd__a22o_1
XFILLER_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$621 U$$621/A _625_/Q VGND VGND VPWR VPWR U$$621/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_37_2 dadda_fa_3_37_2/A dadda_fa_3_37_2/B dadda_fa_3_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/A dadda_fa_4_37_2/B sky130_fd_sc_hd__fa_2
XU$$632 U$$632/A1 U$$682/A2 U$$771/A1 U$$553/X VGND VGND VPWR VPWR U$$633/A sky130_fd_sc_hd__a22o_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$643 U$$643/A U$$661/B VGND VGND VPWR VPWR U$$643/X sky130_fd_sc_hd__xor2_1
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$654 U$$654/A1 U$$682/A2 U$$930/A1 U$$553/X VGND VGND VPWR VPWR U$$655/A sky130_fd_sc_hd__a22o_1
XU$$665 U$$665/A _625_/Q VGND VGND VPWR VPWR U$$665/X sky130_fd_sc_hd__xor2_1
X_585_ _669_/CLK _585_/D VGND VGND VPWR VPWR _585_/Q sky130_fd_sc_hd__dfxtp_4
XU$$676 U$$950/A1 U$$682/A2 U$$952/A1 U$$553/X VGND VGND VPWR VPWR U$$677/A sky130_fd_sc_hd__a22o_1
XU$$687 U$$822/A VGND VGND VPWR VPWR U$$687/Y sky130_fd_sc_hd__inv_1
XFILLER_140_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$698 U$$698/A U$$784/B VGND VGND VPWR VPWR U$$698/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_89_5 dadda_fa_2_89_5/A dadda_fa_2_89_5/B dadda_fa_2_89_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_2/A dadda_fa_4_89_0/A sky130_fd_sc_hd__fa_2
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_26_2 U$$857/X U$$990/X VGND VGND VPWR VPWR dadda_fa_3_27_3/A dadda_fa_4_26_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_32_1 U$$470/X U$$603/X U$$736/X VGND VGND VPWR VPWR dadda_fa_3_33_0/CIN
+ dadda_fa_3_32_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_25_0 U$$57/X U$$190/X U$$323/X VGND VGND VPWR VPWR dadda_fa_3_26_2/CIN
+ dadda_fa_3_25_3/CIN sky130_fd_sc_hd__fa_2
XU$$2050 U$$952/B1 U$$2052/A2 U$$956/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2051/A sky130_fd_sc_hd__a22o_1
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_779__831 VGND VGND VPWR VPWR _779__831/HI U$$4403/B sky130_fd_sc_hd__conb_1
XU$$2061 U$$2061/A1 U$$2059/X _552_/Q U$$2060/X VGND VGND VPWR VPWR U$$2062/A sky130_fd_sc_hd__a22o_1
XU$$2072 U$$2072/A U$$2118/B VGND VGND VPWR VPWR U$$2072/X sky130_fd_sc_hd__xor2_1
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2083 U$$987/A1 U$$2117/A2 U$$28/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2084/A sky130_fd_sc_hd__a22o_1
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2094 U$$2094/A U$$2118/B VGND VGND VPWR VPWR U$$2094/X sky130_fd_sc_hd__xor2_1
XU$$1360 U$$1360/A U$$1369/A VGND VGND VPWR VPWR U$$1360/X sky130_fd_sc_hd__xor2_1
XU$$1371 _636_/Q VGND VGND VPWR VPWR U$$1373/B sky130_fd_sc_hd__inv_1
XU$$1382 U$$971/A1 U$$1474/A2 U$$12/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1383/A sky130_fd_sc_hd__a22o_1
XU$$1393 U$$1393/A U$$1461/B VGND VGND VPWR VPWR U$$1393/X sky130_fd_sc_hd__xor2_1
XFILLER_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_119_1 dadda_fa_5_119_1/A dadda_fa_5_119_1/B dadda_fa_5_119_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_120_0/B dadda_fa_7_119_0/A sky130_fd_sc_hd__fa_1
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_4 U$$2968/X U$$3101/X U$$3234/X VGND VGND VPWR VPWR dadda_fa_2_85_3/B
+ dadda_fa_2_84_5/B sky130_fd_sc_hd__fa_2
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_77_3 U$$2555/X U$$2688/X U$$2821/X VGND VGND VPWR VPWR dadda_fa_2_78_1/B
+ dadda_fa_2_77_4/B sky130_fd_sc_hd__fa_2
XFILLER_131_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_54_2 dadda_fa_4_54_2/A dadda_fa_4_54_2/B dadda_fa_4_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/CIN dadda_fa_5_54_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_47_1 dadda_fa_4_47_1/A dadda_fa_4_47_1/B dadda_fa_4_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/B dadda_fa_5_47_1/B sky130_fd_sc_hd__fa_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_24_0 dadda_fa_7_24_0/A dadda_fa_7_24_0/B dadda_fa_7_24_0/CIN VGND VGND
+ VPWR VPWR _449_/D _320_/D sky130_fd_sc_hd__fa_2
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _499_/CLK _370_/D VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_72_2 U$$1348/X U$$1481/X U$$1614/X VGND VGND VPWR VPWR dadda_fa_1_73_7/CIN
+ dadda_fa_1_72_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_62_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_65_1 U$$536/X U$$669/X U$$802/X VGND VGND VPWR VPWR dadda_fa_1_66_5/CIN
+ dadda_fa_1_65_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_42_0 dadda_fa_3_42_0/A dadda_fa_3_42_0/B dadda_fa_3_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/B dadda_fa_4_42_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_58_0 U$$123/X U$$256/X U$$389/X VGND VGND VPWR VPWR dadda_fa_1_59_6/CIN
+ dadda_fa_1_58_8/A sky130_fd_sc_hd__fa_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$440 U$$440/A U$$530/B VGND VGND VPWR VPWR U$$440/X sky130_fd_sc_hd__xor2_1
X_637_ _637_/CLK _637_/D VGND VGND VPWR VPWR _637_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$451 U$$40/A1 U$$491/A2 _569_/Q U$$416/X VGND VGND VPWR VPWR U$$452/A sky130_fd_sc_hd__a22o_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$462 U$$462/A U$$530/B VGND VGND VPWR VPWR U$$462/X sky130_fd_sc_hd__xor2_1
XFILLER_189_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$473 U$$62/A1 U$$491/A2 U$$64/A1 U$$416/X VGND VGND VPWR VPWR U$$474/A sky130_fd_sc_hd__a22o_1
XU$$484 U$$484/A U$$547/A VGND VGND VPWR VPWR U$$484/X sky130_fd_sc_hd__xor2_1
X_568_ _576_/CLK _568_/D VGND VGND VPWR VPWR _568_/Q sky130_fd_sc_hd__dfxtp_1
XU$$495 U$$84/A1 U$$545/A2 U$$86/A1 U$$416/X VGND VGND VPWR VPWR U$$496/A sky130_fd_sc_hd__a22o_1
XFILLER_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_499_ _499_/CLK _499_/D VGND VGND VPWR VPWR _499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_94_3 U$$3919/X U$$4052/X U$$4185/X VGND VGND VPWR VPWR dadda_fa_3_95_1/B
+ dadda_fa_3_94_3/B sky130_fd_sc_hd__fa_1
XFILLER_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_87_2 U$$4437/X input242/X dadda_fa_2_87_2/CIN VGND VGND VPWR VPWR dadda_fa_3_88_1/A
+ dadda_fa_3_87_3/A sky130_fd_sc_hd__fa_2
XFILLER_113_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_64_1 dadda_fa_5_64_1/A dadda_fa_5_64_1/B dadda_fa_5_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/B dadda_fa_7_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_57_0 dadda_fa_5_57_0/A dadda_fa_5_57_0/B dadda_fa_5_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/A dadda_fa_6_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_8 dadda_fa_1_56_8/A dadda_fa_1_56_8/B dadda_fa_1_56_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_57_3/A dadda_fa_3_56_0/A sky130_fd_sc_hd__fa_2
XFILLER_83_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_103_0 U$$2739/Y U$$2873/X U$$3006/X VGND VGND VPWR VPWR dadda_fa_3_104_2/B
+ dadda_fa_3_103_3/B sky130_fd_sc_hd__fa_2
XFILLER_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1190 U$$92/B1 U$$1218/A2 U$$96/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1191/A sky130_fd_sc_hd__a22o_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_1 U$$1634/X U$$1767/X U$$1900/X VGND VGND VPWR VPWR dadda_fa_2_83_1/CIN
+ dadda_fa_2_82_4/A sky130_fd_sc_hd__fa_2
XFILLER_137_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_75_0 U$$1620/X U$$1753/X U$$1886/X VGND VGND VPWR VPWR dadda_fa_2_76_0/B
+ dadda_fa_2_75_3/B sky130_fd_sc_hd__fa_2
XFILLER_104_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3509 _590_/Q U$$3545/A2 _591_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3510/A sky130_fd_sc_hd__a22o_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2808 U$$4178/A1 U$$2870/A2 _583_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2809/A sky130_fd_sc_hd__a22o_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2819 U$$2819/A U$$2839/B VGND VGND VPWR VPWR U$$2819/X sky130_fd_sc_hd__xor2_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_422_ _645_/CLK _422_/D VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_353_ _490_/CLK _353_/D VGND VGND VPWR VPWR _353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_284_ _612_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_97_1 dadda_fa_3_97_1/A dadda_fa_3_97_1/B dadda_fa_3_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/CIN dadda_fa_4_97_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_74_0 dadda_fa_6_74_0/A dadda_fa_6_74_0/B dadda_fa_6_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_75_0/B dadda_fa_7_74_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_182_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 a[16] VGND VGND VPWR VPWR _632_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_119_0 U$$3835/Y U$$3969/X U$$4102/X VGND VGND VPWR VPWR dadda_fa_5_120_0/CIN
+ dadda_fa_5_119_1/B sky130_fd_sc_hd__fa_2
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$270 U$$270/A _619_/Q VGND VGND VPWR VPWR U$$270/X sky130_fd_sc_hd__xor2_1
XFILLER_189_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$281 U$$281/A U$$357/B VGND VGND VPWR VPWR U$$281/X sky130_fd_sc_hd__xor2_1
XU$$292 U$$975/B1 U$$278/X U$$842/A1 U$$279/X VGND VGND VPWR VPWR U$$293/A sky130_fd_sc_hd__a22o_1
X_741__793 VGND VGND VPWR VPWR _741__793/HI U$$2874/B1 sky130_fd_sc_hd__conb_1
XFILLER_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$6 _430_/Q _302_/Q VGND VGND VPWR VPWR final_adder.U$$6/COUT final_adder.U$$628/A
+ sky130_fd_sc_hd__ha_4
XFILLER_118_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput301 _192_/Q VGND VGND VPWR VPWR o[24] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_0 U$$2984/X U$$3117/X U$$3250/X VGND VGND VPWR VPWR dadda_fa_3_93_0/B
+ dadda_fa_3_92_2/B sky130_fd_sc_hd__fa_2
XFILLER_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput312 _202_/Q VGND VGND VPWR VPWR o[34] sky130_fd_sc_hd__buf_2
Xoutput323 _212_/Q VGND VGND VPWR VPWR o[44] sky130_fd_sc_hd__buf_2
Xoutput334 _222_/Q VGND VGND VPWR VPWR o[54] sky130_fd_sc_hd__buf_2
XFILLER_161_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput345 _232_/Q VGND VGND VPWR VPWR o[64] sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput356 _242_/Q VGND VGND VPWR VPWR o[74] sky130_fd_sc_hd__buf_2
Xoutput367 _252_/Q VGND VGND VPWR VPWR o[84] sky130_fd_sc_hd__buf_2
Xoutput378 _262_/Q VGND VGND VPWR VPWR o[94] sky130_fd_sc_hd__buf_2
XFILLER_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_4_118_2 U$$4499/X input149/X VGND VGND VPWR VPWR dadda_fa_5_119_1/A dadda_ha_4_118_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_114_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_61_6 dadda_fa_1_61_6/A dadda_fa_1_61_6/B dadda_fa_1_61_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/B dadda_fa_2_61_5/B sky130_fd_sc_hd__fa_1
XFILLER_171_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_54_5 U$$2775/X U$$2908/X U$$3041/X VGND VGND VPWR VPWR dadda_fa_2_55_2/A
+ dadda_fa_2_54_5/A sky130_fd_sc_hd__fa_1
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_47_4 U$$1697/X U$$1830/X U$$1963/X VGND VGND VPWR VPWR dadda_fa_2_48_2/CIN
+ dadda_fa_2_47_5/B sky130_fd_sc_hd__fa_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_17_2 dadda_fa_4_17_2/A dadda_fa_4_17_2/B dadda_ha_3_17_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_18_0/CIN dadda_fa_5_17_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_91_0 dadda_fa_7_91_0/A dadda_fa_7_91_0/B dadda_fa_7_91_0/CIN VGND VGND
+ VPWR VPWR _516_/D _387_/D sky130_fd_sc_hd__fa_1
XFILLER_52_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_690__910 VGND VGND VPWR VPWR _690__910/HI _690__910/LO sky130_fd_sc_hd__conb_1
XFILLER_87_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4007 _565_/Q U$$4045/A2 _566_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$4008/A sky130_fd_sc_hd__a22o_1
XU$$4018 U$$4018/A U$$4058/B VGND VGND VPWR VPWR U$$4018/X sky130_fd_sc_hd__xor2_1
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4029 U$$4303/A1 U$$4045/A2 _577_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$4030/A sky130_fd_sc_hd__a22o_1
XFILLER_120_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3306 U$$4265/A1 U$$3396/A2 U$$979/A1 U$$3396/B2 VGND VGND VPWR VPWR U$$3307/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3317 U$$3317/A U$$3397/B VGND VGND VPWR VPWR U$$3317/X sky130_fd_sc_hd__xor2_1
XFILLER_47_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3328 U$$40/A1 U$$3412/A2 U$$3876/B1 U$$3412/B2 VGND VGND VPWR VPWR U$$3329/A sky130_fd_sc_hd__a22o_1
XFILLER_111_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3339 U$$3339/A U$$3397/B VGND VGND VPWR VPWR U$$3339/X sky130_fd_sc_hd__xor2_1
XFILLER_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2605 _655_/Q VGND VGND VPWR VPWR U$$2605/Y sky130_fd_sc_hd__inv_1
XU$$2616 U$$2616/A U$$2710/B VGND VGND VPWR VPWR U$$2616/X sky130_fd_sc_hd__xor2_1
XFILLER_34_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2627 U$$983/A1 U$$2667/A2 U$$4273/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2628/A
+ sky130_fd_sc_hd__a22o_1
XU$$2638 U$$2638/A U$$2694/B VGND VGND VPWR VPWR U$$2638/X sky130_fd_sc_hd__xor2_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_725__777 VGND VGND VPWR VPWR _725__777/HI U$$1915/B1 sky130_fd_sc_hd__conb_1
XU$$2649 U$$4291/B1 U$$2607/X U$$4156/B1 U$$2608/X VGND VGND VPWR VPWR U$$2650/A sky130_fd_sc_hd__a22o_1
XU$$1904 U$$1904/A U$$1904/B VGND VGND VPWR VPWR U$$1904/X sky130_fd_sc_hd__xor2_1
XFILLER_62_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1915 U$$956/A1 U$$1785/X U$$1915/B1 U$$1786/X VGND VGND VPWR VPWR U$$1916/A sky130_fd_sc_hd__a22o_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1926 _552_/Q U$$1922/X U$$969/A1 U$$1923/X VGND VGND VPWR VPWR U$$1927/A sky130_fd_sc_hd__a22o_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1937 U$$1937/A U$$1991/B VGND VGND VPWR VPWR U$$1937/X sky130_fd_sc_hd__xor2_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1948 U$$28/B1 U$$2048/A2 U$$30/B1 U$$2048/B2 VGND VGND VPWR VPWR U$$1949/A sky130_fd_sc_hd__a22o_1
X_405_ _535_/CLK _405_/D VGND VGND VPWR VPWR _405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1959 U$$1959/A U$$1991/B VGND VGND VPWR VPWR U$$1959/X sky130_fd_sc_hd__xor2_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _336_/CLK _336_/D VGND VGND VPWR VPWR _336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_267_ _267_/CLK _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_198_ _329_/CLK _198_/D VGND VGND VPWR VPWR _198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_5 dadda_fa_2_71_5/A dadda_fa_2_71_5/B dadda_fa_2_71_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_2/A dadda_fa_4_71_0/A sky130_fd_sc_hd__fa_2
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_4 dadda_fa_2_64_4/A dadda_fa_2_64_4/B dadda_fa_2_64_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/CIN dadda_fa_3_64_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_57_3 dadda_fa_2_57_3/A dadda_fa_2_57_3/B dadda_fa_2_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/B dadda_fa_3_57_3/B sky130_fd_sc_hd__fa_1
XFILLER_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$11 U$$11/A U$$9/B VGND VGND VPWR VPWR U$$11/X sky130_fd_sc_hd__xor2_1
XU$$22 U$$22/A1 U$$4/X _560_/Q U$$5/X VGND VGND VPWR VPWR U$$23/A sky130_fd_sc_hd__a22o_1
XFILLER_2_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$33 U$$33/A U$$9/B VGND VGND VPWR VPWR U$$33/X sky130_fd_sc_hd__xor2_1
XFILLER_92_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$44 _570_/Q U$$4/X U$$46/A1 U$$5/X VGND VGND VPWR VPWR U$$45/A sky130_fd_sc_hd__a22o_1
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$55 U$$55/A U$$3/A VGND VGND VPWR VPWR U$$55/X sky130_fd_sc_hd__xor2_2
Xdadda_fa_5_27_1 dadda_fa_5_27_1/A dadda_fa_5_27_1/B dadda_fa_5_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/B dadda_fa_7_27_0/A sky130_fd_sc_hd__fa_2
XU$$3840 U$$3838/Y _672_/Q _671_/Q U$$3839/X U$$3836/Y VGND VGND VPWR VPWR U$$3840/X
+ sky130_fd_sc_hd__a32o_4
XU$$66 U$$66/A1 U$$4/X _582_/Q U$$5/X VGND VGND VPWR VPWR U$$67/A sky130_fd_sc_hd__a22o_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3851 U$$3851/A U$$3929/B VGND VGND VPWR VPWR U$$3851/X sky130_fd_sc_hd__xor2_1
XU$$3862 _561_/Q U$$3912/A2 _562_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3863/A sky130_fd_sc_hd__a22o_1
XU$$3873 U$$3873/A U$$3929/B VGND VGND VPWR VPWR U$$3873/X sky130_fd_sc_hd__xor2_1
XU$$77 U$$77/A U$$9/B VGND VGND VPWR VPWR U$$77/X sky130_fd_sc_hd__xor2_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$88 U$$88/A1 U$$4/X U$$90/A1 U$$5/X VGND VGND VPWR VPWR U$$89/A sky130_fd_sc_hd__a22o_1
XU$$3884 U$$4156/B1 U$$3840/X _573_/Q U$$3841/X VGND VGND VPWR VPWR U$$3885/A sky130_fd_sc_hd__a22o_1
XU$$99 U$$99/A U$$3/A VGND VGND VPWR VPWR U$$99/X sky130_fd_sc_hd__xor2_2
XU$$3895 U$$3895/A U$$3929/B VGND VGND VPWR VPWR U$$3895/X sky130_fd_sc_hd__xor2_1
XFILLER_178_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_101_1 dadda_fa_5_101_1/A dadda_fa_5_101_1/B dadda_fa_5_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/B dadda_fa_7_101_0/A sky130_fd_sc_hd__fa_2
XFILLER_174_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_1_39_2 U$$883/X U$$1016/X VGND VGND VPWR VPWR dadda_fa_2_40_4/CIN dadda_fa_3_39_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_52_2 U$$1175/X U$$1308/X U$$1441/X VGND VGND VPWR VPWR dadda_fa_2_53_1/A
+ dadda_fa_2_52_4/A sky130_fd_sc_hd__fa_1
XFILLER_46_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_45_1 U$$496/X U$$629/X U$$762/X VGND VGND VPWR VPWR dadda_fa_2_46_2/B
+ dadda_fa_2_45_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_22_0 dadda_fa_4_22_0/A dadda_fa_4_22_0/B dadda_fa_4_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/A dadda_fa_5_22_1/A sky130_fd_sc_hd__fa_1
XFILLER_44_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_38_0 U$$83/X U$$216/X U$$349/X VGND VGND VPWR VPWR dadda_fa_2_39_4/B dadda_fa_2_38_5/B
+ sky130_fd_sc_hd__fa_2
XFILLER_188_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_74_3 dadda_fa_3_74_3/A dadda_fa_3_74_3/B dadda_fa_3_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/B dadda_fa_4_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_67_2 dadda_fa_3_67_2/A dadda_fa_3_67_2/B dadda_fa_3_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/A dadda_fa_4_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_37_0 dadda_fa_6_37_0/A dadda_fa_6_37_0/B dadda_fa_6_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_38_0/B dadda_fa_7_37_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3103 U$$3103/A U$$3129/B VGND VGND VPWR VPWR U$$3103/X sky130_fd_sc_hd__xor2_1
XU$$3114 _598_/Q U$$3018/X _599_/Q U$$3019/X VGND VGND VPWR VPWR U$$3115/A sky130_fd_sc_hd__a22o_1
XFILLER_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3125 U$$3125/A U$$3137/B VGND VGND VPWR VPWR U$$3125/X sky130_fd_sc_hd__xor2_1
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3136 _609_/Q U$$3018/X _610_/Q U$$3019/X VGND VGND VPWR VPWR U$$3137/A sky130_fd_sc_hd__a22o_1
XU$$2402 U$$2402/A U$$2464/B VGND VGND VPWR VPWR U$$2402/X sky130_fd_sc_hd__xor2_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3147 U$$3147/A _661_/Q VGND VGND VPWR VPWR U$$3147/X sky130_fd_sc_hd__xor2_1
XU$$2413 _590_/Q U$$2421/A2 _591_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2414/A sky130_fd_sc_hd__a22o_1
XU$$3158 U$$3158/A U$$3224/B VGND VGND VPWR VPWR U$$3158/X sky130_fd_sc_hd__xor2_1
XU$$2424 U$$2424/A U$$2436/B VGND VGND VPWR VPWR U$$2424/X sky130_fd_sc_hd__xor2_1
XU$$3169 U$$4265/A1 U$$3243/A2 U$$979/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3170/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2435 U$$928/A1 U$$2463/A2 _602_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2436/A sky130_fd_sc_hd__a22o_1
XFILLER_59_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2446 U$$2446/A U$$2464/B VGND VGND VPWR VPWR U$$2446/X sky130_fd_sc_hd__xor2_1
XU$$1701 U$$1701/A U$$1727/B VGND VGND VPWR VPWR U$$1701/X sky130_fd_sc_hd__xor2_1
XU$$1712 U$$3217/B1 U$$1726/A2 U$$892/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1713/A
+ sky130_fd_sc_hd__a22o_1
XU$$2457 U$$539/A1 U$$2333/X U$$4514/A1 U$$2334/X VGND VGND VPWR VPWR U$$2458/A sky130_fd_sc_hd__a22o_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2468 _653_/Q VGND VGND VPWR VPWR U$$2468/Y sky130_fd_sc_hd__inv_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1723 U$$1723/A U$$1739/B VGND VGND VPWR VPWR U$$1723/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1734 U$$90/A1 U$$1734/A2 U$$92/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1735/A sky130_fd_sc_hd__a22o_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2479 U$$2479/A U$$2533/B VGND VGND VPWR VPWR U$$2479/X sky130_fd_sc_hd__xor2_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1745 U$$1745/A _641_/Q VGND VGND VPWR VPWR U$$1745/X sky130_fd_sc_hd__xor2_1
XU$$1756 _604_/Q U$$1770/A2 U$$799/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1757/A sky130_fd_sc_hd__a22o_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1767 U$$1767/A U$$1781/A VGND VGND VPWR VPWR U$$1767/X sky130_fd_sc_hd__xor2_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1778 U$$956/A1 U$$1648/X U$$1778/B1 U$$1649/X VGND VGND VPWR VPWR U$$1779/A sky130_fd_sc_hd__a22o_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1789 U$$8/A1 U$$1867/A2 U$$8/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1790/A sky130_fd_sc_hd__a22o_1
XFILLER_159_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _452_/CLK _319_/D VGND VGND VPWR VPWR _319_/Q sky130_fd_sc_hd__dfxtp_1
Xinput11 a[19] VGND VGND VPWR VPWR _635_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput22 a[29] VGND VGND VPWR VPWR _645_/D sky130_fd_sc_hd__clkbuf_2
Xinput33 a[39] VGND VGND VPWR VPWR _655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput44 a[49] VGND VGND VPWR VPWR _665_/D sky130_fd_sc_hd__clkbuf_1
Xinput55 a[59] VGND VGND VPWR VPWR _675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput66 b[10] VGND VGND VPWR VPWR _562_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_171_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput77 b[20] VGND VGND VPWR VPWR _572_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_171_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput88 b[30] VGND VGND VPWR VPWR _582_/D sky130_fd_sc_hd__buf_2
Xinput99 b[40] VGND VGND VPWR VPWR _592_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_62_1 dadda_fa_2_62_1/A dadda_fa_2_62_1/B dadda_fa_2_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/CIN dadda_fa_3_62_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater601 _625_/Q VGND VGND VPWR VPWR U$$661/B sky130_fd_sc_hd__buf_12
Xrepeater612 U$$956/A1 VGND VGND VPWR VPWR U$$819/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$419 final_adder.U$$336/B final_adder.U$$686/B final_adder.U$$289/X
+ VGND VGND VPWR VPWR final_adder.U$$690/B sky130_fd_sc_hd__a21o_1
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater623 _610_/Q VGND VGND VPWR VPWR U$$4508/A1 sky130_fd_sc_hd__buf_12
Xrepeater634 U$$4496/A1 VGND VGND VPWR VPWR U$$934/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_55_0 dadda_fa_2_55_0/A dadda_fa_2_55_0/B dadda_fa_2_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/B dadda_fa_3_55_2/B sky130_fd_sc_hd__fa_2
Xrepeater645 _599_/Q VGND VGND VPWR VPWR U$$924/A1 sky130_fd_sc_hd__buf_12
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater656 U$$4476/A1 VGND VGND VPWR VPWR U$$92/A1 sky130_fd_sc_hd__buf_12
Xrepeater667 _590_/Q VGND VGND VPWR VPWR U$$84/A1 sky130_fd_sc_hd__buf_12
XU$$4360 U$$4360/A U$$4384/A VGND VGND VPWR VPWR U$$4360/X sky130_fd_sc_hd__xor2_1
Xrepeater678 U$$76/A1 VGND VGND VPWR VPWR U$$759/B1 sky130_fd_sc_hd__buf_12
XU$$4371 U$$4508/A1 U$$4377/A2 U$$4510/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4372/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater689 U$$3217/B1 VGND VGND VPWR VPWR U$$68/A1 sky130_fd_sc_hd__buf_12
XFILLER_93_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4382 U$$4382/A _679_/Q VGND VGND VPWR VPWR U$$4382/X sky130_fd_sc_hd__xor2_1
XU$$4393 U$$4393/A U$$4393/B VGND VGND VPWR VPWR U$$4393/X sky130_fd_sc_hd__xor2_2
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3670 U$$4492/A1 U$$3566/X U$$4494/A1 U$$3567/X VGND VGND VPWR VPWR U$$3671/A sky130_fd_sc_hd__a22o_1
XU$$3681 U$$3681/A _669_/Q VGND VGND VPWR VPWR U$$3681/X sky130_fd_sc_hd__xor2_1
XFILLER_92_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3692 _613_/Q U$$3566/X U$$4379/A1 U$$3567/X VGND VGND VPWR VPWR U$$3693/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_9_0 U$$291/X U$$424/X U$$557/X VGND VGND VPWR VPWR dadda_fa_6_10_0/A dadda_fa_6_9_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2980 U$$2980/A U$$3004/B VGND VGND VPWR VPWR U$$2980/X sky130_fd_sc_hd__xor2_1
XU$$2991 _605_/Q U$$2881/X _606_/Q U$$2882/X VGND VGND VPWR VPWR U$$2992/A sky130_fd_sc_hd__a22o_1
XFILLER_179_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_84_2 dadda_fa_4_84_2/A dadda_fa_4_84_2/B dadda_fa_4_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/CIN dadda_fa_5_84_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_77_1 dadda_fa_4_77_1/A dadda_fa_4_77_1/B dadda_fa_4_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/B dadda_fa_5_77_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_54_0 dadda_fa_7_54_0/A dadda_fa_7_54_0/B dadda_fa_7_54_0/CIN VGND VGND
+ VPWR VPWR _479_/D _350_/D sky130_fd_sc_hd__fa_1
XFILLER_115_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_670_ _679_/CLK _670_/D VGND VGND VPWR VPWR _670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$803 U$$940/A1 U$$689/X U$$942/A1 U$$690/X VGND VGND VPWR VPWR U$$804/A sky130_fd_sc_hd__a22o_1
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$814 U$$814/A _627_/Q VGND VGND VPWR VPWR U$$814/X sky130_fd_sc_hd__xor2_1
XFILLER_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$825 U$$959/A U$$825/B VGND VGND VPWR VPWR U$$825/X sky130_fd_sc_hd__and2_1
XFILLER_90_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$836 U$$12/B1 U$$928/A2 U$$16/A1 U$$928/B2 VGND VGND VPWR VPWR U$$837/A sky130_fd_sc_hd__a22o_1
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$847 U$$847/A U$$943/B VGND VGND VPWR VPWR U$$847/X sky130_fd_sc_hd__xor2_1
XFILLER_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$858 U$$36/A1 U$$910/A2 U$$38/A1 U$$910/B2 VGND VGND VPWR VPWR U$$859/A sky130_fd_sc_hd__a22o_1
XU$$1008 U$$1008/A U$$992/B VGND VGND VPWR VPWR U$$1008/X sky130_fd_sc_hd__xor2_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$869 U$$869/A U$$903/B VGND VGND VPWR VPWR U$$869/X sky130_fd_sc_hd__xor2_1
XU$$1019 U$$60/A1 U$$963/X U$$62/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1020/A sky130_fd_sc_hd__a22o_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_796__848 VGND VGND VPWR VPWR _796__848/HI U$$4437/B sky130_fd_sc_hd__conb_1
XFILLER_25_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_837__889 VGND VGND VPWR VPWR _837__889/HI U$$5/A2 sky130_fd_sc_hd__conb_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_1_0_1_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_72_0 dadda_fa_3_72_0/A dadda_fa_3_72_0/B dadda_fa_3_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/B dadda_fa_4_72_1/CIN sky130_fd_sc_hd__fa_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2210 U$$18/A1 U$$2196/X U$$20/A1 U$$2197/X VGND VGND VPWR VPWR U$$2211/A sky130_fd_sc_hd__a22o_1
XU$$2221 U$$2221/A U$$2257/B VGND VGND VPWR VPWR U$$2221/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_101_0 dadda_fa_4_101_0/A dadda_fa_4_101_0/B dadda_fa_4_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/A dadda_fa_5_101_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_34_5 U$$2336/X U$$2432/B input184/X VGND VGND VPWR VPWR dadda_fa_3_35_2/A
+ dadda_fa_4_34_0/A sky130_fd_sc_hd__fa_1
XU$$2232 U$$3191/A1 U$$2270/A2 U$$3876/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2233/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2243 U$$2243/A U$$2257/B VGND VGND VPWR VPWR U$$2243/X sky130_fd_sc_hd__xor2_1
XFILLER_23_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2254 U$$3624/A1 U$$2270/A2 U$$3900/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2255/A
+ sky130_fd_sc_hd__a22o_1
XU$$2265 U$$2265/A U$$2327/B VGND VGND VPWR VPWR U$$2265/X sky130_fd_sc_hd__xor2_1
XU$$1520 U$$1520/A U$$1614/B VGND VGND VPWR VPWR U$$1520/X sky130_fd_sc_hd__xor2_1
XU$$2276 _590_/Q U$$2326/A2 _591_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2277/A sky130_fd_sc_hd__a22o_1
XU$$1531 U$$983/A1 U$$1511/X U$$26/A1 U$$1512/X VGND VGND VPWR VPWR U$$1532/A sky130_fd_sc_hd__a22o_1
XU$$1542 U$$1542/A U$$1580/B VGND VGND VPWR VPWR U$$1542/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2287 U$$2287/A U$$2289/B VGND VGND VPWR VPWR U$$2287/X sky130_fd_sc_hd__xor2_1
XU$$1553 U$$46/A1 U$$1511/X _572_/Q U$$1512/X VGND VGND VPWR VPWR U$$1554/A sky130_fd_sc_hd__a22o_1
XU$$2298 _601_/Q U$$2316/A2 U$$928/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2299/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1564 U$$1564/A U$$1580/B VGND VGND VPWR VPWR U$$1564/X sky130_fd_sc_hd__xor2_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1575 U$$3217/B1 U$$1605/A2 U$$892/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1576/A
+ sky130_fd_sc_hd__a22o_1
XU$$1586 U$$1586/A U$$1643/A VGND VGND VPWR VPWR U$$1586/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1597 U$$90/A1 U$$1511/X U$$92/A1 U$$1512/X VGND VGND VPWR VPWR U$$1598/A sky130_fd_sc_hd__a22o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_94_1 dadda_fa_5_94_1/A dadda_fa_5_94_1/B dadda_fa_5_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/B dadda_fa_7_94_0/A sky130_fd_sc_hd__fa_2
XFILLER_163_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_87_0 dadda_fa_5_87_0/A dadda_fa_5_87_0/B dadda_fa_5_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/A dadda_fa_6_87_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_128_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_7 U$$3889/X U$$4022/X U$$4155/X VGND VGND VPWR VPWR dadda_fa_2_80_2/CIN
+ dadda_fa_2_79_5/CIN sky130_fd_sc_hd__fa_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$205 final_adder.U$$699/A final_adder.U$$571/B1 final_adder.U$$205/B1
+ VGND VGND VPWR VPWR final_adder.U$$205/X sky130_fd_sc_hd__a21o_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$216 final_adder.U$$711/A final_adder.U$$710/A VGND VGND VPWR VPWR
+ final_adder.U$$300/B sky130_fd_sc_hd__and2_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater420 U$$2744/X VGND VGND VPWR VPWR U$$2870/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$227 final_adder.U$$721/A final_adder.U$$593/B1 final_adder.U$$227/B1
+ VGND VGND VPWR VPWR final_adder.U$$227/X sky130_fd_sc_hd__a21o_1
Xrepeater431 U$$2059/X VGND VGND VPWR VPWR U$$2117/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$238 final_adder.U$$733/A final_adder.U$$732/A VGND VGND VPWR VPWR
+ final_adder.U$$310/A sky130_fd_sc_hd__and2_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater442 U$$1648/X VGND VGND VPWR VPWR U$$1770/A2 sky130_fd_sc_hd__buf_12
XFILLER_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$249 final_adder.U$$743/A final_adder.U$$615/B1 final_adder.U$$249/B1
+ VGND VGND VPWR VPWR final_adder.U$$249/X sky130_fd_sc_hd__a21o_1
Xrepeater453 U$$964/X VGND VGND VPWR VPWR U$$1073/B2 sky130_fd_sc_hd__buf_12
XFILLER_38_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater464 U$$3978/X VGND VGND VPWR VPWR U$$4063/B2 sky130_fd_sc_hd__buf_12
Xrepeater475 U$$3293/X VGND VGND VPWR VPWR U$$3412/B2 sky130_fd_sc_hd__buf_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater486 U$$2608/X VGND VGND VPWR VPWR U$$2729/B2 sky130_fd_sc_hd__buf_12
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater497 U$$2048/B2 VGND VGND VPWR VPWR U$$2036/B2 sky130_fd_sc_hd__buf_12
XFILLER_53_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4190 U$$765/A1 U$$4114/X _589_/Q U$$4115/X VGND VGND VPWR VPWR U$$4191/A sky130_fd_sc_hd__a22o_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_2 dadda_fa_3_103_2/A dadda_fa_3_103_2/B dadda_fa_3_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/A dadda_fa_4_103_2/B sky130_fd_sc_hd__fa_2
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput201 c[4] VGND VGND VPWR VPWR input201/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput212 c[5] VGND VGND VPWR VPWR input212/X sky130_fd_sc_hd__buf_2
Xinput223 c[6] VGND VGND VPWR VPWR input223/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput234 c[7] VGND VGND VPWR VPWR input234/X sky130_fd_sc_hd__clkbuf_2
Xinput245 c[8] VGND VGND VPWR VPWR input245/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput256 c[9] VGND VGND VPWR VPWR input256/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_67_5 U$$2136/X U$$2269/X U$$2402/X VGND VGND VPWR VPWR dadda_fa_1_68_7/A
+ dadda_fa_2_67_0/A sky130_fd_sc_hd__fa_2
XFILLER_124_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_117_0 dadda_fa_6_117_0/A dadda_fa_6_117_0/B dadda_fa_6_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_118_0/B dadda_fa_7_117_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_653_ _656_/CLK _653_/D VGND VGND VPWR VPWR _653_/Q sky130_fd_sc_hd__dfxtp_4
XU$$600 U$$50/B1 U$$626/A2 U$$876/A1 U$$553/X VGND VGND VPWR VPWR U$$601/A sky130_fd_sc_hd__a22o_1
XU$$611 U$$611/A U$$661/B VGND VGND VPWR VPWR U$$611/X sky130_fd_sc_hd__xor2_1
XU$$622 U$$759/A1 U$$626/A2 U$$759/B1 U$$553/X VGND VGND VPWR VPWR U$$623/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_37_3 dadda_fa_3_37_3/A dadda_fa_3_37_3/B dadda_fa_3_37_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/B dadda_fa_4_37_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$633 U$$633/A _625_/Q VGND VGND VPWR VPWR U$$633/X sky130_fd_sc_hd__xor2_1
XU$$644 U$$96/A1 U$$682/A2 U$$96/B1 U$$553/X VGND VGND VPWR VPWR U$$645/A sky130_fd_sc_hd__a22o_1
XU$$655 U$$655/A _625_/Q VGND VGND VPWR VPWR U$$655/X sky130_fd_sc_hd__xor2_1
X_584_ _594_/CLK _584_/D VGND VGND VPWR VPWR _584_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$666 U$$940/A1 U$$552/X U$$942/A1 U$$553/X VGND VGND VPWR VPWR U$$667/A sky130_fd_sc_hd__a22o_1
XU$$677 U$$677/A _625_/Q VGND VGND VPWR VPWR U$$677/X sky130_fd_sc_hd__xor2_1
XU$$688 U$$822/A U$$688/B VGND VGND VPWR VPWR U$$688/X sky130_fd_sc_hd__and2_1
XFILLER_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$699 U$$12/B1 U$$817/A2 U$$16/A1 U$$785/B2 VGND VGND VPWR VPWR U$$700/A sky130_fd_sc_hd__a22o_1
XFILLER_140_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_32_2 U$$869/X U$$1002/X U$$1135/X VGND VGND VPWR VPWR dadda_fa_3_33_1/A
+ dadda_fa_3_32_3/A sky130_fd_sc_hd__fa_2
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2040 U$$944/A1 U$$2052/A2 U$$946/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2041/A sky130_fd_sc_hd__a22o_1
XU$$2051 U$$2051/A U$$2055/A VGND VGND VPWR VPWR U$$2051/X sky130_fd_sc_hd__xor2_1
XU$$2062 U$$2062/A U$$2186/B VGND VGND VPWR VPWR U$$2062/X sky130_fd_sc_hd__xor2_1
XU$$2073 U$$4265/A1 U$$2117/A2 U$$979/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2074/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2084 U$$2084/A U$$2118/B VGND VGND VPWR VPWR U$$2084/X sky130_fd_sc_hd__xor2_1
XU$$1350 U$$1350/A _635_/Q VGND VGND VPWR VPWR U$$1350/X sky130_fd_sc_hd__xor2_1
XU$$2095 U$$3191/A1 U$$2117/A2 U$$3876/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2096/A
+ sky130_fd_sc_hd__a22o_1
XU$$1361 U$$539/A1 U$$1367/A2 U$$4514/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1362/A
+ sky130_fd_sc_hd__a22o_1
XU$$1372 _637_/Q VGND VGND VPWR VPWR U$$1372/Y sky130_fd_sc_hd__inv_1
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1383 U$$1383/A U$$1479/B VGND VGND VPWR VPWR U$$1383/X sky130_fd_sc_hd__xor2_1
XU$$1394 _560_/Q U$$1474/A2 U$$26/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1395/A sky130_fd_sc_hd__a22o_1
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_84_5 U$$3367/X U$$3500/X U$$3633/X VGND VGND VPWR VPWR dadda_fa_2_85_3/CIN
+ dadda_fa_2_84_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_77_4 U$$2954/X U$$3087/X U$$3220/X VGND VGND VPWR VPWR dadda_fa_2_78_1/CIN
+ dadda_fa_2_77_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_47_2 dadda_fa_4_47_2/A dadda_fa_4_47_2/B dadda_fa_4_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/CIN dadda_fa_5_47_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_17_0 dadda_fa_7_17_0/A dadda_fa_7_17_0/B dadda_fa_7_17_0/CIN VGND VGND
+ VPWR VPWR _442_/D _313_/D sky130_fd_sc_hd__fa_2
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$90 _514_/Q _386_/Q VGND VGND VPWR VPWR final_adder.U$$585/B1 final_adder.U$$712/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_59_3 U$$1322/X U$$1455/X VGND VGND VPWR VPWR dadda_fa_1_60_7/B dadda_fa_2_59_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_150_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_65_2 U$$935/X U$$1068/X U$$1201/X VGND VGND VPWR VPWR dadda_fa_1_66_6/A
+ dadda_fa_1_65_8/A sky130_fd_sc_hd__fa_1
XFILLER_97_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_42_1 dadda_fa_3_42_1/A dadda_fa_3_42_1/B dadda_fa_3_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/CIN dadda_fa_4_42_2/A sky130_fd_sc_hd__fa_2
Xdadda_fa_0_58_1 U$$522/X U$$655/X U$$788/X VGND VGND VPWR VPWR dadda_fa_1_59_7/A
+ dadda_fa_1_58_8/B sky130_fd_sc_hd__fa_2
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_35_0 dadda_fa_3_35_0/A dadda_fa_3_35_0/B dadda_fa_3_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/B dadda_fa_4_35_1/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$591 final_adder.U$$718/A final_adder.U$$718/B final_adder.U$$591/B1
+ VGND VGND VPWR VPWR final_adder.U$$719/B sky130_fd_sc_hd__a21o_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$430 U$$430/A U$$547/A VGND VGND VPWR VPWR U$$430/X sky130_fd_sc_hd__xor2_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$441 U$$28/B1 U$$491/A2 U$$32/A1 U$$416/X VGND VGND VPWR VPWR U$$442/A sky130_fd_sc_hd__a22o_1
X_636_ _642_/CLK _636_/D VGND VGND VPWR VPWR _636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$452 U$$452/A U$$530/B VGND VGND VPWR VPWR U$$452/X sky130_fd_sc_hd__xor2_1
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$463 U$$52/A1 U$$545/A2 U$$54/A1 U$$416/X VGND VGND VPWR VPWR U$$464/A sky130_fd_sc_hd__a22o_1
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$474 U$$474/A U$$547/A VGND VGND VPWR VPWR U$$474/X sky130_fd_sc_hd__xor2_1
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$485 U$$759/A1 U$$491/A2 U$$759/B1 U$$416/X VGND VGND VPWR VPWR U$$486/A sky130_fd_sc_hd__a22o_1
X_567_ _637_/CLK _567_/D VGND VGND VPWR VPWR _567_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$496 U$$496/A U$$547/A VGND VGND VPWR VPWR U$$496/X sky130_fd_sc_hd__xor2_1
XFILLER_60_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_498_ _501_/CLK _498_/D VGND VGND VPWR VPWR _498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_94_4 U$$4318/X U$$4451/X input250/X VGND VGND VPWR VPWR dadda_fa_3_95_1/CIN
+ dadda_fa_3_94_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_87_3 dadda_fa_2_87_3/A dadda_fa_2_87_3/B dadda_fa_2_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/B dadda_fa_3_87_3/B sky130_fd_sc_hd__fa_1
XFILLER_153_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_57_1 dadda_fa_5_57_1/A dadda_fa_5_57_1/B dadda_fa_5_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/B dadda_fa_7_57_0/A sky130_fd_sc_hd__fa_1
XFILLER_80_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_103_1 U$$3139/X U$$3272/X U$$3405/X VGND VGND VPWR VPWR dadda_fa_3_104_2/CIN
+ dadda_fa_3_103_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1180 U$$84/A1 U$$1218/A2 U$$908/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1181/A sky130_fd_sc_hd__a22o_1
XU$$1191 U$$1191/A U$$1232/A VGND VGND VPWR VPWR U$$1191/X sky130_fd_sc_hd__xor2_1
XFILLER_176_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_124_0 _703__923/HI U$$4245/X U$$4378/X VGND VGND VPWR VPWR dadda_fa_6_125_0/B
+ dadda_fa_6_124_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_149_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_82_2 U$$2033/X U$$2166/X U$$2299/X VGND VGND VPWR VPWR dadda_fa_2_83_2/A
+ dadda_fa_2_82_4/B sky130_fd_sc_hd__fa_1
XFILLER_131_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_75_1 U$$2019/X U$$2152/X U$$2285/X VGND VGND VPWR VPWR dadda_fa_2_76_0/CIN
+ dadda_fa_2_75_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_52_0 dadda_fa_4_52_0/A dadda_fa_4_52_0/B dadda_fa_4_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/A dadda_fa_5_52_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_68_0 U$$2537/X U$$2670/X U$$2803/X VGND VGND VPWR VPWR dadda_fa_2_69_0/B
+ dadda_fa_2_68_3/B sky130_fd_sc_hd__fa_2
Xdadda_ha_2_102_3 U$$3802/X U$$3935/X VGND VGND VPWR VPWR dadda_fa_3_103_3/A dadda_fa_4_102_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_86_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2809 U$$2809/A U$$2839/B VGND VGND VPWR VPWR U$$2809/X sky130_fd_sc_hd__xor2_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_421_ _677_/CLK _421_/D VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_clk _560_/CLK VGND VGND VPWR VPWR _639_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _483_/CLK _352_/D VGND VGND VPWR VPWR _352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_283_ _612_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_97_2 dadda_fa_3_97_2/A dadda_fa_3_97_2/B dadda_fa_3_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/A dadda_fa_4_97_2/B sky130_fd_sc_hd__fa_2
XFILLER_142_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_67_0 dadda_fa_6_67_0/A dadda_fa_6_67_0/B dadda_fa_6_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_68_0/B dadda_fa_7_67_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_70_0 _681__901/HI U$$546/X U$$679/X VGND VGND VPWR VPWR dadda_fa_1_71_6/B
+ dadda_fa_1_70_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 a[17] VGND VGND VPWR VPWR _633_/D sky130_fd_sc_hd__buf_2
XFILLER_188_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_119_1 U$$4235/X U$$4368/X U$$4501/X VGND VGND VPWR VPWR dadda_fa_5_120_1/A
+ dadda_fa_5_119_1/CIN sky130_fd_sc_hd__fa_2
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_5_6_1 U$$418/X U$$547/A VGND VGND VPWR VPWR dadda_fa_6_7_0/B dadda_fa_7_6_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$260 U$$260/A U$$262/B VGND VGND VPWR VPWR U$$260/X sky130_fd_sc_hd__xor2_1
XFILLER_18_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$271 U$$819/A1 U$$141/X U$$271/B1 U$$142/X VGND VGND VPWR VPWR U$$272/A sky130_fd_sc_hd__a22o_1
XFILLER_33_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_619_ _642_/CLK _619_/D VGND VGND VPWR VPWR _619_/Q sky130_fd_sc_hd__dfxtp_4
XU$$282 U$$8/A1 U$$278/X U$$8/B1 U$$279/X VGND VGND VPWR VPWR U$$283/A sky130_fd_sc_hd__a22o_1
XFILLER_189_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$293 U$$293/A U$$391/B VGND VGND VPWR VPWR U$$293/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_71_clk _560_/CLK VGND VGND VPWR VPWR _669_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$7 _431_/Q _303_/Q VGND VGND VPWR VPWR final_adder.U$$7/COUT final_adder.U$$7/SUM
+ sky130_fd_sc_hd__ha_4
Xoutput302 _193_/Q VGND VGND VPWR VPWR o[25] sky130_fd_sc_hd__buf_2
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_92_1 U$$3383/X U$$3516/X U$$3649/X VGND VGND VPWR VPWR dadda_fa_3_93_0/CIN
+ dadda_fa_3_92_2/CIN sky130_fd_sc_hd__fa_2
Xoutput313 _203_/Q VGND VGND VPWR VPWR o[35] sky130_fd_sc_hd__buf_2
Xoutput324 _213_/Q VGND VGND VPWR VPWR o[45] sky130_fd_sc_hd__buf_2
Xoutput335 _223_/Q VGND VGND VPWR VPWR o[55] sky130_fd_sc_hd__buf_2
Xoutput346 _233_/Q VGND VGND VPWR VPWR o[65] sky130_fd_sc_hd__buf_2
XFILLER_142_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_85_0 U$$3901/X U$$4034/X U$$4167/X VGND VGND VPWR VPWR dadda_fa_3_86_0/B
+ dadda_fa_3_85_2/B sky130_fd_sc_hd__fa_2
XFILLER_160_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput357 _243_/Q VGND VGND VPWR VPWR o[75] sky130_fd_sc_hd__buf_2
Xoutput368 _253_/Q VGND VGND VPWR VPWR o[85] sky130_fd_sc_hd__buf_2
Xoutput379 _263_/Q VGND VGND VPWR VPWR o[95] sky130_fd_sc_hd__buf_2
XFILLER_87_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_48_7 U$$2896/X U$$3029/X VGND VGND VPWR VPWR dadda_fa_2_49_3/B dadda_fa_3_48_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_61_7 dadda_fa_1_61_7/A dadda_fa_1_61_7/B dadda_fa_1_61_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/CIN dadda_fa_2_61_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_54_6 U$$3174/X U$$3307/X U$$3440/X VGND VGND VPWR VPWR dadda_fa_2_55_2/B
+ dadda_fa_2_54_5/B sky130_fd_sc_hd__fa_1
XFILLER_110_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_47_5 U$$2096/X U$$2229/X U$$2362/X VGND VGND VPWR VPWR dadda_fa_2_48_3/A
+ dadda_fa_2_47_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_167_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_6_0 dadda_fa_7_6_0/A dadda_fa_7_6_0/B dadda_fa_7_6_0/CIN VGND VGND VPWR
+ VPWR _431_/D _302_/D sky130_fd_sc_hd__fa_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_62_clk _536_/CLK VGND VGND VPWR VPWR _583_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_84_0 dadda_fa_7_84_0/A dadda_fa_7_84_0/B dadda_fa_7_84_0/CIN VGND VGND
+ VPWR VPWR _509_/D _380_/D sky130_fd_sc_hd__fa_2
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4008 U$$4008/A U$$4044/B VGND VGND VPWR VPWR U$$4008/X sky130_fd_sc_hd__xor2_1
XU$$4019 U$$4291/B1 U$$3977/X U$$4156/B1 U$$3978/X VGND VGND VPWR VPWR U$$4020/A sky130_fd_sc_hd__a22o_1
XFILLER_150_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3307 U$$3307/A U$$3397/B VGND VGND VPWR VPWR U$$3307/X sky130_fd_sc_hd__xor2_1
XU$$3318 U$$30/A1 U$$3396/A2 U$$30/B1 U$$3396/B2 VGND VGND VPWR VPWR U$$3319/A sky130_fd_sc_hd__a22o_1
XU$$3329 U$$3329/A U$$3413/B VGND VGND VPWR VPWR U$$3329/X sky130_fd_sc_hd__xor2_1
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2606 _655_/Q U$$2606/B VGND VGND VPWR VPWR U$$2606/X sky130_fd_sc_hd__and2_1
XFILLER_111_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2617 U$$14/A1 U$$2667/A2 U$$14/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2618/A sky130_fd_sc_hd__a22o_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2628 U$$2628/A U$$2694/B VGND VGND VPWR VPWR U$$2628/X sky130_fd_sc_hd__xor2_1
XU$$2639 U$$4283/A1 U$$2667/A2 U$$4285/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2640/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1905 U$$4508/A1 U$$1785/X U$$4510/A1 U$$1786/X VGND VGND VPWR VPWR U$$1906/A sky130_fd_sc_hd__a22o_1
XFILLER_15_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1916 U$$1916/A _643_/Q VGND VGND VPWR VPWR U$$1916/X sky130_fd_sc_hd__xor2_2
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1927 U$$1927/A U$$2021/B VGND VGND VPWR VPWR U$$1927/X sky130_fd_sc_hd__xor2_2
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1938 U$$979/A1 U$$2036/A2 U$$979/B1 U$$2036/B2 VGND VGND VPWR VPWR U$$1939/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_53_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _518_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_404_ _535_/CLK _404_/D VGND VGND VPWR VPWR _404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1949 U$$1949/A U$$1991/B VGND VGND VPWR VPWR U$$1949/X sky130_fd_sc_hd__xor2_1
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _463_/CLK _335_/D VGND VGND VPWR VPWR _335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_266_ _280_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_197_ _329_/CLK _197_/D VGND VGND VPWR VPWR _197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_64_5 dadda_fa_2_64_5/A dadda_fa_2_64_5/B dadda_fa_2_64_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_2/A dadda_fa_4_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_57_4 dadda_fa_2_57_4/A dadda_fa_2_57_4/B dadda_fa_2_57_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/CIN dadda_fa_3_57_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_65_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$12 U$$12/A1 U$$4/X U$$12/B1 U$$5/X VGND VGND VPWR VPWR U$$13/A sky130_fd_sc_hd__a22o_1
XU$$23 U$$23/A U$$89/B VGND VGND VPWR VPWR U$$23/X sky130_fd_sc_hd__xor2_1
XU$$34 U$$34/A1 U$$4/X U$$36/A1 U$$5/X VGND VGND VPWR VPWR U$$35/A sky130_fd_sc_hd__a22o_1
XU$$3830 U$$3830/A U$$3835/A VGND VGND VPWR VPWR U$$3830/X sky130_fd_sc_hd__xor2_1
XU$$45 U$$45/A U$$3/A VGND VGND VPWR VPWR U$$45/X sky130_fd_sc_hd__xor2_1
XFILLER_92_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3841 U$$3839/B _671_/Q _672_/Q U$$3836/Y VGND VGND VPWR VPWR U$$3841/X sky130_fd_sc_hd__a22o_4
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$56 U$$56/A1 U$$4/X U$$58/A1 U$$5/X VGND VGND VPWR VPWR U$$57/A sky130_fd_sc_hd__a22o_1
XU$$67 U$$67/A U$$89/B VGND VGND VPWR VPWR U$$67/X sky130_fd_sc_hd__xor2_2
XU$$3852 _556_/Q U$$3840/X U$$975/B1 U$$3841/X VGND VGND VPWR VPWR U$$3853/A sky130_fd_sc_hd__a22o_1
XU$$78 U$$78/A1 U$$4/X U$$80/A1 U$$5/X VGND VGND VPWR VPWR U$$79/A sky130_fd_sc_hd__a22o_1
XU$$3863 U$$3863/A U$$3893/B VGND VGND VPWR VPWR U$$3863/X sky130_fd_sc_hd__xor2_1
XU$$3874 U$$4285/A1 U$$3840/X U$$4424/A1 U$$3841/X VGND VGND VPWR VPWR U$$3875/A sky130_fd_sc_hd__a22o_1
XU$$3885 U$$3885/A U$$3929/B VGND VGND VPWR VPWR U$$3885/X sky130_fd_sc_hd__xor2_1
XU$$89 U$$89/A U$$89/B VGND VGND VPWR VPWR U$$89/X sky130_fd_sc_hd__xor2_1
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3896 U$$4170/A1 U$$3912/A2 U$$4446/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3897/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_44_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _267_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_52_3 U$$1574/X U$$1707/X U$$1840/X VGND VGND VPWR VPWR dadda_fa_2_53_1/B
+ dadda_fa_2_52_4/B sky130_fd_sc_hd__fa_1
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_45_2 U$$895/X U$$1028/X U$$1161/X VGND VGND VPWR VPWR dadda_fa_2_46_2/CIN
+ dadda_fa_2_45_5/A sky130_fd_sc_hd__fa_2
XFILLER_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_22_1 dadda_fa_4_22_1/A dadda_fa_4_22_1/B dadda_fa_4_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/B dadda_fa_5_22_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_38_1 U$$482/X U$$615/X U$$748/X VGND VGND VPWR VPWR dadda_fa_2_39_4/CIN
+ dadda_fa_2_38_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_35_clk _369_/CLK VGND VGND VPWR VPWR _496_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_4_15_0 U$$303/X U$$436/X U$$569/X VGND VGND VPWR VPWR dadda_fa_5_16_0/A
+ dadda_fa_5_15_1/A sky130_fd_sc_hd__fa_1
XFILLER_24_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_67_3 dadda_fa_3_67_3/A dadda_fa_3_67_3/B dadda_fa_3_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/B dadda_fa_4_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3104 U$$912/A1 U$$3146/A2 U$$4476/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3105/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3115 U$$3115/A U$$3137/B VGND VGND VPWR VPWR U$$3115/X sky130_fd_sc_hd__xor2_1
XFILLER_19_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3126 _604_/Q U$$3018/X _605_/Q U$$3019/X VGND VGND VPWR VPWR U$$3127/A sky130_fd_sc_hd__a22o_1
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3137 U$$3137/A U$$3137/B VGND VGND VPWR VPWR U$$3137/X sky130_fd_sc_hd__xor2_1
XU$$3148 U$$819/A1 U$$3018/X U$$3148/B1 U$$3019/X VGND VGND VPWR VPWR U$$3149/A sky130_fd_sc_hd__a22o_1
XU$$2403 U$$74/A1 U$$2421/A2 U$$2953/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2404/A sky130_fd_sc_hd__a22o_1
XU$$2414 U$$2414/A U$$2436/B VGND VGND VPWR VPWR U$$2414/X sky130_fd_sc_hd__xor2_1
XFILLER_34_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3159 U$$8/A1 U$$3241/A2 U$$969/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3160/A sky130_fd_sc_hd__a22o_1
XFILLER_59_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2425 U$$96/A1 U$$2463/A2 _597_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2426/A sky130_fd_sc_hd__a22o_1
XU$$2436 U$$2436/A U$$2436/B VGND VGND VPWR VPWR U$$2436/X sky130_fd_sc_hd__xor2_1
XU$$1702 U$$58/A1 U$$1734/A2 U$$60/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1703/A sky130_fd_sc_hd__a22o_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2447 _607_/Q U$$2463/A2 _608_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2448/A sky130_fd_sc_hd__a22o_1
XU$$1713 U$$1713/A U$$1739/B VGND VGND VPWR VPWR U$$1713/X sky130_fd_sc_hd__xor2_1
XFILLER_27_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2458 U$$2458/A U$$2464/B VGND VGND VPWR VPWR U$$2458/X sky130_fd_sc_hd__xor2_1
XFILLER_188_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_clk _369_/CLK VGND VGND VPWR VPWR _483_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1724 U$$80/A1 U$$1734/A2 U$$82/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1725/A sky130_fd_sc_hd__a22o_1
XU$$2469 _653_/Q U$$2469/B VGND VGND VPWR VPWR U$$2469/X sky130_fd_sc_hd__and2_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1735 U$$1735/A U$$1781/A VGND VGND VPWR VPWR U$$1735/X sky130_fd_sc_hd__xor2_1
X_697__917 VGND VGND VPWR VPWR _697__917/HI _697__917/LO sky130_fd_sc_hd__conb_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1746 _599_/Q U$$1770/A2 _600_/Q U$$1770/B2 VGND VGND VPWR VPWR U$$1747/A sky130_fd_sc_hd__a22o_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1757 U$$1757/A _641_/Q VGND VGND VPWR VPWR U$$1757/X sky130_fd_sc_hd__xor2_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1768 _610_/Q U$$1770/A2 _611_/Q U$$1770/B2 VGND VGND VPWR VPWR U$$1769/A sky130_fd_sc_hd__a22o_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1779 U$$1779/A U$$1781/A VGND VGND VPWR VPWR U$$1779/X sky130_fd_sc_hd__xor2_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_318_ _452_/CLK _318_/D VGND VGND VPWR VPWR _318_/Q sky130_fd_sc_hd__dfxtp_1
Xinput12 a[1] VGND VGND VPWR VPWR _617_/D sky130_fd_sc_hd__buf_4
XFILLER_168_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput23 a[2] VGND VGND VPWR VPWR _618_/D sky130_fd_sc_hd__buf_6
Xinput34 a[3] VGND VGND VPWR VPWR _619_/D sky130_fd_sc_hd__clkbuf_4
X_249_ _379_/CLK _249_/D VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_1
Xinput45 a[4] VGND VGND VPWR VPWR _620_/D sky130_fd_sc_hd__buf_6
XFILLER_156_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput56 a[5] VGND VGND VPWR VPWR _621_/D sky130_fd_sc_hd__buf_4
Xinput67 b[11] VGND VGND VPWR VPWR _563_/D sky130_fd_sc_hd__clkbuf_4
Xinput78 b[21] VGND VGND VPWR VPWR _573_/D sky130_fd_sc_hd__clkbuf_4
Xinput89 b[31] VGND VGND VPWR VPWR _583_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_170_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_62_2 dadda_fa_2_62_2/A dadda_fa_2_62_2/B dadda_fa_2_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/A dadda_fa_3_62_3/A sky130_fd_sc_hd__fa_2
Xrepeater602 _623_/Q VGND VGND VPWR VPWR U$$530/B sky130_fd_sc_hd__buf_12
XFILLER_112_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$409 final_adder.U$$326/B final_adder.U$$646/B final_adder.U$$269/X
+ VGND VGND VPWR VPWR final_adder.U$$650/B sky130_fd_sc_hd__a21o_1
Xrepeater613 _615_/Q VGND VGND VPWR VPWR U$$956/A1 sky130_fd_sc_hd__buf_12
Xrepeater624 U$$4506/A1 VGND VGND VPWR VPWR U$$944/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_55_1 dadda_fa_2_55_1/A dadda_fa_2_55_1/B dadda_fa_2_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/CIN dadda_fa_3_55_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_111_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater635 _604_/Q VGND VGND VPWR VPWR U$$4496/A1 sky130_fd_sc_hd__buf_12
Xrepeater646 _599_/Q VGND VGND VPWR VPWR U$$4486/A1 sky130_fd_sc_hd__buf_12
Xrepeater657 U$$4476/A1 VGND VGND VPWR VPWR U$$914/A1 sky130_fd_sc_hd__buf_12
XU$$4350 U$$4350/A _679_/Q VGND VGND VPWR VPWR U$$4350/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_32_0 dadda_fa_5_32_0/A dadda_fa_5_32_0/B dadda_fa_5_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/A dadda_fa_6_32_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater668 _590_/Q VGND VGND VPWR VPWR U$$632/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_48_0 U$$3162/X U$$3295/X U$$3413/B VGND VGND VPWR VPWR dadda_fa_3_49_0/B
+ dadda_fa_3_48_2/B sky130_fd_sc_hd__fa_2
Xrepeater679 _586_/Q VGND VGND VPWR VPWR U$$76/A1 sky130_fd_sc_hd__buf_12
XU$$4361 U$$936/A1 U$$4377/A2 U$$4500/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4362/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4372 U$$4372/A U$$4384/A VGND VGND VPWR VPWR U$$4372/X sky130_fd_sc_hd__xor2_1
XU$$4383 U$$4384/A VGND VGND VPWR VPWR U$$4383/Y sky130_fd_sc_hd__inv_1
XFILLER_93_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4394 _553_/Q U$$4388/X _554_/Q U$$4389/X VGND VGND VPWR VPWR U$$4395/A sky130_fd_sc_hd__a22o_1
XFILLER_19_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3660 U$$98/A1 U$$3678/A2 U$$98/B1 U$$3678/B2 VGND VGND VPWR VPWR U$$3661/A sky130_fd_sc_hd__a22o_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3671 U$$3671/A U$$3698/A VGND VGND VPWR VPWR U$$3671/X sky130_fd_sc_hd__xor2_1
XFILLER_53_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3682 U$$4504/A1 U$$3566/X U$$4506/A1 U$$3567/X VGND VGND VPWR VPWR U$$3683/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _452_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3693 U$$3693/A U$$3698/A VGND VGND VPWR VPWR U$$3693/X sky130_fd_sc_hd__xor2_1
XFILLER_179_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2970 U$$2970/A _659_/Q VGND VGND VPWR VPWR U$$2970/X sky130_fd_sc_hd__xor2_1
XFILLER_178_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2981 _600_/Q U$$2881/X _601_/Q U$$2882/X VGND VGND VPWR VPWR U$$2982/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_9_1 input256/X dadda_fa_5_9_1/B dadda_ha_4_9_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_6_10_0/B dadda_fa_7_9_0/A sky130_fd_sc_hd__fa_2
XU$$2992 U$$2992/A U$$3004/B VGND VGND VPWR VPWR U$$2992/X sky130_fd_sc_hd__xor2_1
XFILLER_61_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_77_2 dadda_fa_4_77_2/A dadda_fa_4_77_2/B dadda_fa_4_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/CIN dadda_fa_5_77_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_47_0 dadda_fa_7_47_0/A dadda_fa_7_47_0/B dadda_fa_7_47_0/CIN VGND VGND
+ VPWR VPWR _472_/D _343_/D sky130_fd_sc_hd__fa_2
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_50_0 U$$107/X U$$240/X U$$373/X VGND VGND VPWR VPWR dadda_fa_2_51_0/B
+ dadda_fa_2_50_3/B sky130_fd_sc_hd__fa_2
XU$$804 U$$804/A U$$822/A VGND VGND VPWR VPWR U$$804/X sky130_fd_sc_hd__xor2_1
XU$$815 U$$952/A1 U$$817/A2 U$$952/B1 U$$817/B2 VGND VGND VPWR VPWR U$$816/A sky130_fd_sc_hd__a22o_1
XU$$826 U$$824/Y _628_/Q U$$822/A U$$825/X U$$822/Y VGND VGND VPWR VPWR U$$826/X sky130_fd_sc_hd__a32o_4
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$837 U$$837/A U$$959/A VGND VGND VPWR VPWR U$$837/X sky130_fd_sc_hd__xor2_1
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$848 U$$26/A1 U$$928/A2 U$$987/A1 U$$928/B2 VGND VGND VPWR VPWR U$$849/A sky130_fd_sc_hd__a22o_1
XFILLER_83_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$859 U$$859/A U$$923/B VGND VGND VPWR VPWR U$$859/X sky130_fd_sc_hd__xor2_1
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1009 U$$50/A1 U$$999/A2 U$$2790/B1 U$$987/B2 VGND VGND VPWR VPWR U$$1010/A sky130_fd_sc_hd__a22o_1
XFILLER_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_72_1 dadda_fa_3_72_1/A dadda_fa_3_72_1/B dadda_fa_3_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/CIN dadda_fa_4_72_2/A sky130_fd_sc_hd__fa_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_65_0 dadda_fa_3_65_0/A dadda_fa_3_65_0/B dadda_fa_3_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/B dadda_fa_4_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2200 U$$8/A1 U$$2270/A2 U$$8/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2201/A sky130_fd_sc_hd__a22o_1
XFILLER_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2211 U$$2211/A U$$2289/B VGND VGND VPWR VPWR U$$2211/X sky130_fd_sc_hd__xor2_1
XFILLER_35_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_101_1 dadda_fa_4_101_1/A dadda_fa_4_101_1/B dadda_fa_4_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/B dadda_fa_5_101_1/B sky130_fd_sc_hd__fa_1
XU$$2222 U$$30/A1 U$$2270/A2 U$$30/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2223/A sky130_fd_sc_hd__a22o_1
XFILLER_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2233 U$$2233/A U$$2257/B VGND VGND VPWR VPWR U$$2233/X sky130_fd_sc_hd__xor2_1
XU$$2244 U$$2790/B1 U$$2270/A2 U$$4438/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2245/A
+ sky130_fd_sc_hd__a22o_1
XU$$1510 _639_/Q U$$1510/B VGND VGND VPWR VPWR U$$1510/X sky130_fd_sc_hd__and2_1
XU$$2255 U$$2255/A U$$2289/B VGND VGND VPWR VPWR U$$2255/X sky130_fd_sc_hd__xor2_1
XFILLER_179_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1521 U$$12/B1 U$$1511/X U$$16/A1 U$$1512/X VGND VGND VPWR VPWR U$$1522/A sky130_fd_sc_hd__a22o_1
XFILLER_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2266 U$$759/A1 U$$2196/X U$$759/B1 U$$2197/X VGND VGND VPWR VPWR U$$2267/A sky130_fd_sc_hd__a22o_1
XFILLER_50_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2277 U$$2277/A U$$2289/B VGND VGND VPWR VPWR U$$2277/X sky130_fd_sc_hd__xor2_1
XU$$1532 U$$1532/A U$$1614/B VGND VGND VPWR VPWR U$$1532/X sky130_fd_sc_hd__xor2_1
XU$$2288 _596_/Q U$$2326/A2 _597_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2289/A sky130_fd_sc_hd__a22o_1
X_820__872 VGND VGND VPWR VPWR _820__872/HI U$$4485/B sky130_fd_sc_hd__conb_1
XU$$1543 U$$36/A1 U$$1511/X U$$38/A1 U$$1512/X VGND VGND VPWR VPWR U$$1544/A sky130_fd_sc_hd__a22o_1
XFILLER_188_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1554 U$$1554/A U$$1614/B VGND VGND VPWR VPWR U$$1554/X sky130_fd_sc_hd__xor2_1
XU$$2299 U$$2299/A U$$2327/B VGND VGND VPWR VPWR U$$2299/X sky130_fd_sc_hd__xor2_1
XU$$1565 U$$58/A1 U$$1591/A2 U$$60/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1566/A sky130_fd_sc_hd__a22o_1
XFILLER_188_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1576 U$$1576/A U$$1580/B VGND VGND VPWR VPWR U$$1576/X sky130_fd_sc_hd__xor2_1
XFILLER_188_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1587 _588_/Q U$$1641/A2 U$$902/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1588/A sky130_fd_sc_hd__a22o_1
XFILLER_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_122_0 dadda_fa_7_122_0/A dadda_fa_7_122_0/B dadda_fa_7_122_0/CIN VGND
+ VGND VPWR VPWR _547_/D _418_/D sky130_fd_sc_hd__fa_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1598 U$$1598/A _639_/Q VGND VGND VPWR VPWR U$$1598/X sky130_fd_sc_hd__xor2_1
XFILLER_179_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_87_1 dadda_fa_5_87_1/A dadda_fa_5_87_1/B dadda_fa_5_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/B dadda_fa_7_87_0/A sky130_fd_sc_hd__fa_2
XFILLER_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_6_clk _431_/CLK VGND VGND VPWR VPWR _467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_8 U$$4288/X U$$4421/X input233/X VGND VGND VPWR VPWR dadda_fa_2_80_3/A
+ dadda_fa_3_79_0/A sky130_fd_sc_hd__fa_2
XFILLER_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$206 final_adder.U$$701/A final_adder.U$$700/A VGND VGND VPWR VPWR
+ final_adder.U$$294/A sky130_fd_sc_hd__and2_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater410 U$$3292/X VGND VGND VPWR VPWR U$$3396/A2 sky130_fd_sc_hd__buf_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$217 final_adder.U$$711/A final_adder.U$$583/B1 final_adder.U$$217/B1
+ VGND VGND VPWR VPWR final_adder.U$$217/X sky130_fd_sc_hd__a21o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater421 U$$2729/A2 VGND VGND VPWR VPWR U$$2667/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$228 final_adder.U$$723/A final_adder.U$$722/A VGND VGND VPWR VPWR
+ final_adder.U$$306/B sky130_fd_sc_hd__and2_1
Xrepeater432 U$$2189/A2 VGND VGND VPWR VPWR U$$2161/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$239 final_adder.U$$733/A final_adder.U$$605/B1 final_adder.U$$239/B1
+ VGND VGND VPWR VPWR final_adder.U$$239/X sky130_fd_sc_hd__a21o_1
Xrepeater443 U$$1591/A2 VGND VGND VPWR VPWR U$$1605/A2 sky130_fd_sc_hd__buf_12
Xrepeater454 U$$964/X VGND VGND VPWR VPWR U$$999/B2 sky130_fd_sc_hd__buf_12
XFILLER_73_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater465 U$$3841/X VGND VGND VPWR VPWR U$$3912/B2 sky130_fd_sc_hd__buf_12
Xrepeater476 U$$3156/X VGND VGND VPWR VPWR U$$3243/B2 sky130_fd_sc_hd__buf_12
XFILLER_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater487 U$$2584/B2 VGND VGND VPWR VPWR U$$2534/B2 sky130_fd_sc_hd__buf_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater498 U$$2052/B2 VGND VGND VPWR VPWR U$$2048/B2 sky130_fd_sc_hd__buf_12
XU$$4180 U$$70/A1 U$$4244/A2 U$$70/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4181/A sky130_fd_sc_hd__a22o_1
XFILLER_38_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4191 U$$4191/A U$$4247/A VGND VGND VPWR VPWR U$$4191/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3490 U$$3490/A _667_/Q VGND VGND VPWR VPWR U$$3490/X sky130_fd_sc_hd__xor2_1
XFILLER_43_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_82_0 dadda_fa_4_82_0/A dadda_fa_4_82_0/B dadda_fa_4_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/A dadda_fa_5_82_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_3 dadda_fa_3_103_3/A dadda_fa_3_103_3/B dadda_fa_3_103_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/B dadda_fa_4_103_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput202 c[50] VGND VGND VPWR VPWR input202/X sky130_fd_sc_hd__buf_4
Xinput213 c[60] VGND VGND VPWR VPWR input213/X sky130_fd_sc_hd__clkbuf_2
Xinput224 c[70] VGND VGND VPWR VPWR input224/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput235 c[80] VGND VGND VPWR VPWR input235/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput246 c[90] VGND VGND VPWR VPWR input246/X sky130_fd_sc_hd__buf_2
X_763__815 VGND VGND VPWR VPWR _763__815/HI U$$417/A1 sky130_fd_sc_hd__conb_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$740 final_adder.U$$740/A final_adder.U$$740/B VGND VGND VPWR VPWR
+ _286_/D sky130_fd_sc_hd__xor2_1
XFILLER_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_652_ _667_/CLK _652_/D VGND VGND VPWR VPWR _652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$601 U$$601/A U$$623/B VGND VGND VPWR VPWR U$$601/X sky130_fd_sc_hd__xor2_1
XU$$612 U$$64/A1 U$$682/A2 U$$66/A1 U$$553/X VGND VGND VPWR VPWR U$$613/A sky130_fd_sc_hd__a22o_1
XU$$623 U$$623/A U$$623/B VGND VGND VPWR VPWR U$$623/X sky130_fd_sc_hd__xor2_1
XU$$634 U$$86/A1 U$$682/A2 U$$88/A1 U$$553/X VGND VGND VPWR VPWR U$$635/A sky130_fd_sc_hd__a22o_1
XFILLER_90_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$645 U$$645/A U$$661/B VGND VGND VPWR VPWR U$$645/X sky130_fd_sc_hd__xor2_1
X_804__856 VGND VGND VPWR VPWR _804__856/HI U$$4453/B sky130_fd_sc_hd__conb_1
XFILLER_90_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_583_ _583_/CLK _583_/D VGND VGND VPWR VPWR _583_/Q sky130_fd_sc_hd__dfxtp_4
XU$$656 U$$930/A1 U$$682/A2 U$$932/A1 U$$553/X VGND VGND VPWR VPWR U$$657/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$667 U$$667/A _625_/Q VGND VGND VPWR VPWR U$$667/X sky130_fd_sc_hd__xor2_1
XFILLER_44_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$678 U$$952/A1 U$$682/A2 U$$952/B1 U$$553/X VGND VGND VPWR VPWR U$$679/A sky130_fd_sc_hd__a22o_1
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$689 U$$687/Y _626_/Q _625_/Q U$$688/X U$$685/Y VGND VGND VPWR VPWR U$$689/X sky130_fd_sc_hd__a32o_4
XFILLER_44_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_97_0 dadda_fa_6_97_0/A dadda_fa_6_97_0/B dadda_fa_6_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_98_0/B dadda_fa_7_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_8_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_2_33_5 U$$2068/X U$$2201/X VGND VGND VPWR VPWR dadda_fa_3_34_2/A dadda_fa_4_33_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_32_3 U$$1268/X U$$1401/X U$$1534/X VGND VGND VPWR VPWR dadda_fa_3_33_1/B
+ dadda_fa_3_32_3/B sky130_fd_sc_hd__fa_2
XU$$2030 U$$4496/A1 U$$2048/A2 U$$799/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$2031/A
+ sky130_fd_sc_hd__a22o_1
XU$$2041 U$$2041/A U$$2055/A VGND VGND VPWR VPWR U$$2041/X sky130_fd_sc_hd__xor2_1
XU$$2052 U$$956/A1 U$$2052/A2 U$$2052/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2053/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2063 _552_/Q U$$2059/X U$$969/A1 U$$2060/X VGND VGND VPWR VPWR U$$2064/A sky130_fd_sc_hd__a22o_1
XU$$2074 U$$2074/A U$$2118/B VGND VGND VPWR VPWR U$$2074/X sky130_fd_sc_hd__xor2_1
XFILLER_35_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1340 U$$1340/A U$$1369/A VGND VGND VPWR VPWR U$$1340/X sky130_fd_sc_hd__xor2_1
XU$$2085 U$$28/B1 U$$2117/A2 U$$30/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2086/A sky130_fd_sc_hd__a22o_1
XFILLER_16_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2096 U$$2096/A U$$2118/B VGND VGND VPWR VPWR U$$2096/X sky130_fd_sc_hd__xor2_1
XU$$1351 _607_/Q U$$1367/A2 _608_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1352/A sky130_fd_sc_hd__a22o_1
XU$$1362 U$$1362/A _635_/Q VGND VGND VPWR VPWR U$$1362/X sky130_fd_sc_hd__xor2_1
XU$$1373 _637_/Q U$$1373/B VGND VGND VPWR VPWR U$$1373/X sky130_fd_sc_hd__and2_1
XFILLER_148_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1384 U$$14/A1 U$$1474/A2 U$$14/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1385/A sky130_fd_sc_hd__a22o_1
XU$$1395 U$$1395/A U$$1479/B VGND VGND VPWR VPWR U$$1395/X sky130_fd_sc_hd__xor2_1
XFILLER_188_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_77_5 U$$3353/X U$$3486/X U$$3619/X VGND VGND VPWR VPWR dadda_fa_2_78_2/A
+ dadda_fa_2_77_5/A sky130_fd_sc_hd__fa_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$80 _504_/Q _376_/Q VGND VGND VPWR VPWR final_adder.U$$575/B1 final_adder.U$$702/A
+ sky130_fd_sc_hd__ha_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$91 _515_/Q _387_/Q VGND VGND VPWR VPWR final_adder.U$$219/B1 final_adder.U$$713/A
+ sky130_fd_sc_hd__ha_2
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_101_0 U$$4199/X U$$4332/X U$$4465/X VGND VGND VPWR VPWR dadda_fa_4_102_0/B
+ dadda_fa_4_101_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_65_3 U$$1334/X U$$1467/X U$$1600/X VGND VGND VPWR VPWR dadda_fa_1_66_6/B
+ dadda_fa_1_65_8/B sky130_fd_sc_hd__fa_1
XFILLER_130_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_42_2 dadda_fa_3_42_2/A dadda_fa_3_42_2/B dadda_fa_3_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/A dadda_fa_4_42_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_58_2 U$$921/X U$$1054/X U$$1187/X VGND VGND VPWR VPWR dadda_fa_1_59_7/B
+ dadda_fa_1_58_8/CIN sky130_fd_sc_hd__fa_2
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_35_1 dadda_fa_3_35_1/A dadda_fa_3_35_1/B dadda_fa_3_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/CIN dadda_fa_4_35_2/A sky130_fd_sc_hd__fa_2
XFILLER_57_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$581 final_adder.U$$708/A final_adder.U$$708/B final_adder.U$$581/B1
+ VGND VGND VPWR VPWR final_adder.U$$709/B sky130_fd_sc_hd__a21o_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$420 U$$420/A U$$530/B VGND VGND VPWR VPWR U$$420/X sky130_fd_sc_hd__xor2_1
X_635_ _646_/CLK _635_/D VGND VGND VPWR VPWR _635_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$431 U$$20/A1 U$$491/A2 _559_/Q U$$416/X VGND VGND VPWR VPWR U$$432/A sky130_fd_sc_hd__a22o_1
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$442 U$$442/A U$$530/B VGND VGND VPWR VPWR U$$442/X sky130_fd_sc_hd__xor2_1
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$453 _569_/Q U$$491/A2 _570_/Q U$$416/X VGND VGND VPWR VPWR U$$454/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_12_0 dadda_fa_6_12_0/A dadda_fa_6_12_0/B dadda_fa_6_12_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_13_0/B dadda_fa_7_12_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_91_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$464 U$$464/A U$$530/B VGND VGND VPWR VPWR U$$464/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_28_0 U$$1526/X U$$1659/X U$$1792/X VGND VGND VPWR VPWR dadda_fa_4_29_0/B
+ dadda_fa_4_28_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_566_ _576_/CLK _566_/D VGND VGND VPWR VPWR _566_/Q sky130_fd_sc_hd__dfxtp_4
XU$$475 U$$64/A1 U$$491/A2 U$$66/A1 U$$416/X VGND VGND VPWR VPWR U$$476/A sky130_fd_sc_hd__a22o_1
XU$$486 U$$486/A U$$530/B VGND VGND VPWR VPWR U$$486/X sky130_fd_sc_hd__xor2_1
XFILLER_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$497 U$$86/A1 U$$545/A2 U$$88/A1 U$$416/X VGND VGND VPWR VPWR U$$498/A sky130_fd_sc_hd__a22o_1
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_497_ _497_/CLK _497_/D VGND VGND VPWR VPWR _497_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_160_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_94_5 dadda_fa_2_94_5/A dadda_fa_2_94_5/B dadda_fa_2_94_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_95_2/A dadda_fa_4_94_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_87_4 dadda_fa_2_87_4/A dadda_fa_2_87_4/B dadda_fa_2_87_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/CIN dadda_fa_3_87_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_24_1 U$$454/X U$$587/X VGND VGND VPWR VPWR dadda_fa_3_25_3/B dadda_fa_4_24_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_30_0 U$$67/X U$$200/X U$$333/X VGND VGND VPWR VPWR dadda_fa_3_31_1/A dadda_fa_3_30_2/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_165_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_103_2 U$$3538/X U$$3671/X U$$3804/X VGND VGND VPWR VPWR dadda_fa_3_104_3/A
+ dadda_fa_4_103_0/A sky130_fd_sc_hd__fa_2
XFILLER_39_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1170 U$$759/A1 U$$1200/A2 U$$759/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1171/A sky130_fd_sc_hd__a22o_1
XU$$1181 U$$1181/A U$$1232/A VGND VGND VPWR VPWR U$$1181/X sky130_fd_sc_hd__xor2_1
XU$$1192 U$$96/A1 U$$1218/A2 U$$96/B1 U$$1218/B2 VGND VGND VPWR VPWR U$$1193/A sky130_fd_sc_hd__a22o_1
XFILLER_188_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_117_0 dadda_fa_5_117_0/A dadda_fa_5_117_0/B dadda_fa_5_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/A dadda_fa_6_117_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_3 U$$2432/X U$$2565/X U$$2698/X VGND VGND VPWR VPWR dadda_fa_2_83_2/B
+ dadda_fa_2_82_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_75_2 U$$2418/X U$$2551/X U$$2684/X VGND VGND VPWR VPWR dadda_fa_2_76_1/A
+ dadda_fa_2_75_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_52_1 dadda_fa_4_52_1/A dadda_fa_4_52_1/B dadda_fa_4_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/B dadda_fa_5_52_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_68_1 U$$2936/X U$$3069/X U$$3202/X VGND VGND VPWR VPWR dadda_fa_2_69_0/CIN
+ dadda_fa_2_68_3/CIN sky130_fd_sc_hd__fa_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_45_0 dadda_fa_4_45_0/A dadda_fa_4_45_0/B dadda_fa_4_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/A dadda_fa_5_45_1/A sky130_fd_sc_hd__fa_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_420_ _656_/CLK _420_/D VGND VGND VPWR VPWR _420_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_351_ _480_/CLK _351_/D VGND VGND VPWR VPWR _351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_282_ _612_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_97_3 dadda_fa_3_97_3/A dadda_fa_3_97_3/B dadda_fa_3_97_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/B dadda_fa_4_97_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_182_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_769__821 VGND VGND VPWR VPWR _769__821/HI U$$4387/A sky130_fd_sc_hd__conb_1
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_70_1 U$$812/X U$$945/X U$$1078/X VGND VGND VPWR VPWR dadda_fa_1_71_6/CIN
+ dadda_fa_1_70_8/A sky130_fd_sc_hd__fa_2
XFILLER_104_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_63_0 U$$133/X U$$266/X U$$399/X VGND VGND VPWR VPWR dadda_fa_1_64_5/B
+ dadda_fa_1_63_7/B sky130_fd_sc_hd__fa_2
XFILLER_76_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$250 U$$250/A U$$274/A VGND VGND VPWR VPWR U$$250/X sky130_fd_sc_hd__xor2_1
X_618_ _620_/CLK _618_/D VGND VGND VPWR VPWR _618_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$261 U$$946/A1 U$$141/X U$$948/A1 U$$142/X VGND VGND VPWR VPWR U$$262/A sky130_fd_sc_hd__a22o_1
XFILLER_91_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$272 U$$272/A _619_/Q VGND VGND VPWR VPWR U$$272/X sky130_fd_sc_hd__xor2_1
XFILLER_33_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$283 U$$283/A U$$357/B VGND VGND VPWR VPWR U$$283/X sky130_fd_sc_hd__xor2_1
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$294 U$$842/A1 U$$278/X U$$22/A1 U$$279/X VGND VGND VPWR VPWR U$$295/A sky130_fd_sc_hd__a22o_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ _594_/CLK _549_/D VGND VGND VPWR VPWR _549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$0 U$$0/A VGND VGND VPWR VPWR U$$0/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$8 _432_/Q _304_/Q VGND VGND VPWR VPWR final_adder.U$$8/COUT final_adder.U$$8/SUM
+ sky130_fd_sc_hd__ha_2
XFILLER_133_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput303 _194_/Q VGND VGND VPWR VPWR o[26] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_2 U$$3782/X U$$3915/X U$$4048/X VGND VGND VPWR VPWR dadda_fa_3_93_1/A
+ dadda_fa_3_92_3/A sky130_fd_sc_hd__fa_1
Xoutput314 _204_/Q VGND VGND VPWR VPWR o[36] sky130_fd_sc_hd__buf_2
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput325 _214_/Q VGND VGND VPWR VPWR o[46] sky130_fd_sc_hd__buf_2
Xoutput336 _224_/Q VGND VGND VPWR VPWR o[56] sky130_fd_sc_hd__buf_2
Xoutput347 _234_/Q VGND VGND VPWR VPWR o[66] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_1 U$$4300/X U$$4433/X input240/X VGND VGND VPWR VPWR dadda_fa_3_86_0/CIN
+ dadda_fa_3_85_2/CIN sky130_fd_sc_hd__fa_2
Xoutput358 _244_/Q VGND VGND VPWR VPWR o[76] sky130_fd_sc_hd__buf_2
Xoutput369 _254_/Q VGND VGND VPWR VPWR o[86] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_62_0 dadda_fa_5_62_0/A dadda_fa_5_62_0/B dadda_fa_5_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/A dadda_fa_6_62_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_78_0 dadda_fa_2_78_0/A dadda_fa_2_78_0/B dadda_fa_2_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/B dadda_fa_3_78_2/B sky130_fd_sc_hd__fa_2
XFILLER_113_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_61_8 dadda_fa_1_61_8/A dadda_fa_1_61_8/B dadda_fa_1_61_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_3/A dadda_fa_3_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_54_7 U$$3573/X U$$3706/X U$$3756/B VGND VGND VPWR VPWR dadda_fa_2_55_2/CIN
+ dadda_fa_2_54_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_77_0 dadda_fa_7_77_0/A dadda_fa_7_77_0/B dadda_fa_7_77_0/CIN VGND VGND
+ VPWR VPWR _502_/D _373_/D sky130_fd_sc_hd__fa_1
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_80_0 _685__905/HI U$$1231/X U$$1364/X VGND VGND VPWR VPWR dadda_fa_2_81_0/CIN
+ dadda_fa_2_80_3/B sky130_fd_sc_hd__fa_1
XFILLER_133_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4009 _566_/Q U$$4045/A2 _567_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$4010/A sky130_fd_sc_hd__a22o_1
XFILLER_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3308 U$$842/A1 U$$3412/A2 U$$22/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3309/A sky130_fd_sc_hd__a22o_1
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3319 U$$3319/A U$$3397/B VGND VGND VPWR VPWR U$$3319/X sky130_fd_sc_hd__xor2_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2607 U$$2605/Y _654_/Q U$$2603/A U$$2606/X U$$2603/Y VGND VGND VPWR VPWR U$$2607/X
+ sky130_fd_sc_hd__a32o_4
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2618 U$$2618/A U$$2694/B VGND VGND VPWR VPWR U$$2618/X sky130_fd_sc_hd__xor2_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2629 _561_/Q U$$2667/A2 U$$28/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2630/A sky130_fd_sc_hd__a22o_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1906 U$$1906/A _643_/Q VGND VGND VPWR VPWR U$$1906/X sky130_fd_sc_hd__xor2_1
XFILLER_55_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1917 _643_/Q VGND VGND VPWR VPWR U$$1917/Y sky130_fd_sc_hd__inv_1
XU$$1928 U$$969/A1 U$$1922/X U$$12/A1 U$$1923/X VGND VGND VPWR VPWR U$$1929/A sky130_fd_sc_hd__a22o_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1939 U$$1939/A U$$1991/B VGND VGND VPWR VPWR U$$1939/X sky130_fd_sc_hd__xor2_1
XFILLER_26_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _537_/CLK _403_/D VGND VGND VPWR VPWR _403_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _448_/CLK _334_/D VGND VGND VPWR VPWR _334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_265_ _267_/CLK _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_196_ _333_/CLK _196_/D VGND VGND VPWR VPWR _196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_95_0 dadda_fa_3_95_0/A dadda_fa_3_95_0/B dadda_fa_3_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/B dadda_fa_4_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4510 U$$4510/A1 U$$4388/X U$$539/A1 U$$4389/X VGND VGND VPWR VPWR U$$4511/A sky130_fd_sc_hd__a22o_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_57_5 dadda_fa_2_57_5/A dadda_fa_2_57_5/B dadda_fa_2_57_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_2/A dadda_fa_4_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_38_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$13 U$$13/A U$$9/B VGND VGND VPWR VPWR U$$13/X sky130_fd_sc_hd__xor2_1
XU$$24 _560_/Q U$$4/X U$$26/A1 U$$5/X VGND VGND VPWR VPWR U$$25/A sky130_fd_sc_hd__a22o_1
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$35 U$$35/A U$$3/A VGND VGND VPWR VPWR U$$35/X sky130_fd_sc_hd__xor2_1
XU$$3820 U$$3820/A U$$3835/A VGND VGND VPWR VPWR U$$3820/X sky130_fd_sc_hd__xor2_1
XFILLER_65_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3831 U$$4379/A1 U$$3703/X U$$819/A1 U$$3704/X VGND VGND VPWR VPWR U$$3832/A sky130_fd_sc_hd__a22o_1
XU$$46 U$$46/A1 U$$4/X _572_/Q U$$5/X VGND VGND VPWR VPWR U$$47/A sky130_fd_sc_hd__a22o_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3842 U$$3842/A1 U$$3912/A2 U$$4255/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3843/A
+ sky130_fd_sc_hd__a22o_1
XU$$57 U$$57/A U$$3/A VGND VGND VPWR VPWR U$$57/X sky130_fd_sc_hd__xor2_1
XFILLER_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3853 U$$3853/A U$$3929/B VGND VGND VPWR VPWR U$$3853/X sky130_fd_sc_hd__xor2_1
XU$$68 U$$68/A1 U$$4/X U$$68/B1 U$$5/X VGND VGND VPWR VPWR U$$69/A sky130_fd_sc_hd__a22o_1
XU$$3864 _562_/Q U$$3912/A2 _563_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3865/A sky130_fd_sc_hd__a22o_1
XU$$79 U$$79/A U$$3/A VGND VGND VPWR VPWR U$$79/X sky130_fd_sc_hd__xor2_1
XFILLER_46_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3875 U$$3875/A U$$3929/B VGND VGND VPWR VPWR U$$3875/X sky130_fd_sc_hd__xor2_1
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3886 _573_/Q U$$3840/X _574_/Q U$$3841/X VGND VGND VPWR VPWR U$$3887/A sky130_fd_sc_hd__a22o_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3897 U$$3897/A U$$3929/B VGND VGND VPWR VPWR U$$3897/X sky130_fd_sc_hd__xor2_1
XFILLER_45_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_4 U$$1973/X U$$2106/X U$$2239/X VGND VGND VPWR VPWR dadda_fa_2_53_1/CIN
+ dadda_fa_2_52_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_45_3 U$$1294/X U$$1427/X U$$1560/X VGND VGND VPWR VPWR dadda_fa_2_46_3/A
+ dadda_fa_2_45_5/B sky130_fd_sc_hd__fa_2
XFILLER_56_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_22_2 dadda_fa_4_22_2/A dadda_fa_4_22_2/B dadda_fa_4_22_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/CIN dadda_fa_5_22_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_15_1 U$$702/X U$$835/X U$$968/X VGND VGND VPWR VPWR dadda_fa_5_16_0/B
+ dadda_fa_5_15_1/B sky130_fd_sc_hd__fa_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_731__783 VGND VGND VPWR VPWR _731__783/HI U$$2326/B1 sky130_fd_sc_hd__conb_1
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3105 U$$3105/A U$$3129/B VGND VGND VPWR VPWR U$$3105/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3116 _599_/Q U$$3018/X _600_/Q U$$3019/X VGND VGND VPWR VPWR U$$3117/A sky130_fd_sc_hd__a22o_1
XU$$3127 U$$3127/A U$$3137/B VGND VGND VPWR VPWR U$$3127/X sky130_fd_sc_hd__xor2_1
XU$$3138 U$$4508/A1 U$$3146/A2 U$$4510/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3139/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2404 U$$2404/A U$$2432/B VGND VGND VPWR VPWR U$$2404/X sky130_fd_sc_hd__xor2_1
XFILLER_35_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3149 U$$3149/A _661_/Q VGND VGND VPWR VPWR U$$3149/X sky130_fd_sc_hd__xor2_1
XU$$2415 _591_/Q U$$2463/A2 U$$4335/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2416/A sky130_fd_sc_hd__a22o_1
XFILLER_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2426 U$$2426/A U$$2464/B VGND VGND VPWR VPWR U$$2426/X sky130_fd_sc_hd__xor2_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2437 U$$4492/A1 U$$2463/A2 U$$4494/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2438/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1703 U$$1703/A U$$1781/A VGND VGND VPWR VPWR U$$1703/X sky130_fd_sc_hd__xor2_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2448 U$$2448/A U$$2464/B VGND VGND VPWR VPWR U$$2448/X sky130_fd_sc_hd__xor2_1
XU$$1714 U$$892/A1 U$$1726/A2 U$$892/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1715/A sky130_fd_sc_hd__a22o_1
XU$$2459 _613_/Q U$$2463/A2 _614_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2460/A sky130_fd_sc_hd__a22o_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1725 U$$1725/A U$$1781/A VGND VGND VPWR VPWR U$$1725/X sky130_fd_sc_hd__xor2_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1736 U$$92/A1 U$$1770/A2 U$$92/B1 U$$1770/B2 VGND VGND VPWR VPWR U$$1737/A sky130_fd_sc_hd__a22o_1
XU$$1747 U$$1747/A _641_/Q VGND VGND VPWR VPWR U$$1747/X sky130_fd_sc_hd__xor2_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1758 U$$799/A1 U$$1648/X U$$938/A1 U$$1649/X VGND VGND VPWR VPWR U$$1759/A sky130_fd_sc_hd__a22o_1
XU$$1769 U$$1769/A _641_/Q VGND VGND VPWR VPWR U$$1769/X sky130_fd_sc_hd__xor2_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_317_ _452_/CLK _317_/D VGND VGND VPWR VPWR _317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput13 a[20] VGND VGND VPWR VPWR _636_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_248_ _267_/CLK _248_/D VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput24 a[30] VGND VGND VPWR VPWR _646_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 a[40] VGND VGND VPWR VPWR _656_/D sky130_fd_sc_hd__clkbuf_1
Xinput46 a[50] VGND VGND VPWR VPWR _666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput57 a[60] VGND VGND VPWR VPWR _676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput68 b[12] VGND VGND VPWR VPWR _564_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_179_ _336_/CLK _179_/D VGND VGND VPWR VPWR _179_/Q sky130_fd_sc_hd__dfxtp_1
Xinput79 b[22] VGND VGND VPWR VPWR _574_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_62_3 dadda_fa_2_62_3/A dadda_fa_2_62_3/B dadda_fa_2_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/B dadda_fa_3_62_3/B sky130_fd_sc_hd__fa_1
Xrepeater603 _623_/Q VGND VGND VPWR VPWR U$$547/A sky130_fd_sc_hd__buf_12
XFILLER_42_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater614 U$$4379/A1 VGND VGND VPWR VPWR U$$952/B1 sky130_fd_sc_hd__buf_12
XFILLER_42_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater625 _609_/Q VGND VGND VPWR VPWR U$$4506/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_55_2 dadda_fa_2_55_2/A dadda_fa_2_55_2/B dadda_fa_2_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/A dadda_fa_3_55_3/A sky130_fd_sc_hd__fa_1
XFILLER_84_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater636 U$$4494/A1 VGND VGND VPWR VPWR U$$932/A1 sky130_fd_sc_hd__buf_12
Xrepeater647 U$$4484/A1 VGND VGND VPWR VPWR U$$98/B1 sky130_fd_sc_hd__buf_12
XFILLER_111_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater658 _594_/Q VGND VGND VPWR VPWR U$$4476/A1 sky130_fd_sc_hd__buf_12
X_680__900 VGND VGND VPWR VPWR _680__900/HI _680__900/LO sky130_fd_sc_hd__conb_1
XU$$4340 U$$4340/A _679_/Q VGND VGND VPWR VPWR U$$4340/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_32_1 dadda_fa_5_32_1/A dadda_fa_5_32_1/B dadda_fa_5_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/B dadda_fa_7_32_0/A sky130_fd_sc_hd__fa_1
Xrepeater669 _589_/Q VGND VGND VPWR VPWR U$$902/B1 sky130_fd_sc_hd__buf_12
XU$$4351 U$$787/B1 U$$4377/A2 U$$654/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4352/A sky130_fd_sc_hd__a22o_1
XU$$4362 U$$4362/A U$$4384/A VGND VGND VPWR VPWR U$$4362/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_1 input199/X dadda_fa_2_48_1/B dadda_fa_2_48_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_49_0/CIN dadda_fa_3_48_2/CIN sky130_fd_sc_hd__fa_2
XU$$4373 U$$4510/A1 U$$4377/A2 U$$539/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4374/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4384 U$$4384/A VGND VGND VPWR VPWR U$$4384/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_5_25_0 dadda_fa_5_25_0/A dadda_fa_5_25_0/B dadda_fa_5_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/A dadda_fa_6_25_0/CIN sky130_fd_sc_hd__fa_1
XU$$4395 U$$4395/A U$$4395/B VGND VGND VPWR VPWR U$$4395/X sky130_fd_sc_hd__xor2_2
XU$$3650 U$$771/B1 U$$3678/A2 U$$90/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3651/A sky130_fd_sc_hd__a22o_1
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3661 U$$3661/A _669_/Q VGND VGND VPWR VPWR U$$3661/X sky130_fd_sc_hd__xor2_1
XFILLER_19_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3672 U$$4494/A1 U$$3678/A2 U$$934/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3673/A
+ sky130_fd_sc_hd__a22o_1
XU$$3683 U$$3683/A U$$3698/A VGND VGND VPWR VPWR U$$3683/X sky130_fd_sc_hd__xor2_1
XFILLER_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3694 U$$4379/A1 U$$3566/X U$$819/A1 U$$3567/X VGND VGND VPWR VPWR U$$3695/A sky130_fd_sc_hd__a22o_1
XU$$2960 U$$2960/A U$$2960/B VGND VGND VPWR VPWR U$$2960/X sky130_fd_sc_hd__xor2_1
XU$$2971 U$$92/B1 U$$2975/A2 U$$96/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2972/A sky130_fd_sc_hd__a22o_1
XU$$2982 U$$2982/A U$$3004/B VGND VGND VPWR VPWR U$$2982/X sky130_fd_sc_hd__xor2_1
XU$$2993 _606_/Q U$$3009/A2 U$$940/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2994/A sky130_fd_sc_hd__a22o_1
XFILLER_179_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_715__767 VGND VGND VPWR VPWR _715__767/HI U$$134/B1 sky130_fd_sc_hd__conb_1
XFILLER_173_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_1_37_1 U$$480/X U$$613/X VGND VGND VPWR VPWR dadda_fa_2_38_5/A dadda_fa_3_37_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_29_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_50_1 U$$506/X U$$639/X U$$772/X VGND VGND VPWR VPWR dadda_fa_2_51_0/CIN
+ dadda_fa_2_50_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_84_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$805 U$$942/A1 U$$689/X U$$944/A1 U$$690/X VGND VGND VPWR VPWR U$$806/A sky130_fd_sc_hd__a22o_1
XFILLER_56_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$816 U$$816/A _627_/Q VGND VGND VPWR VPWR U$$816/X sky130_fd_sc_hd__xor2_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$827 U$$825/B U$$822/A _628_/Q U$$822/Y VGND VGND VPWR VPWR U$$827/X sky130_fd_sc_hd__a22o_4
Xdadda_fa_1_43_0 U$$93/X U$$226/X U$$359/X VGND VGND VPWR VPWR dadda_fa_2_44_2/CIN
+ dadda_fa_2_43_4/CIN sky130_fd_sc_hd__fa_1
XU$$838 U$$16/A1 U$$928/A2 U$$975/B1 U$$928/B2 VGND VGND VPWR VPWR U$$839/A sky130_fd_sc_hd__a22o_1
XU$$849 U$$849/A U$$923/B VGND VGND VPWR VPWR U$$849/X sky130_fd_sc_hd__xor2_1
XFILLER_71_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_72_2 dadda_fa_3_72_2/A dadda_fa_3_72_2/B dadda_fa_3_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/A dadda_fa_4_72_2/B sky130_fd_sc_hd__fa_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_65_1 dadda_fa_3_65_1/A dadda_fa_3_65_1/B dadda_fa_3_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/CIN dadda_fa_4_65_2/A sky130_fd_sc_hd__fa_1
XFILLER_154_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_42_0 dadda_fa_6_42_0/A dadda_fa_6_42_0/B dadda_fa_6_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_43_0/B dadda_fa_7_42_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_58_0 dadda_fa_3_58_0/A dadda_fa_3_58_0/B dadda_fa_3_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/B dadda_fa_4_58_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2201 U$$2201/A U$$2257/B VGND VGND VPWR VPWR U$$2201/X sky130_fd_sc_hd__xor2_1
X_705__925 VGND VGND VPWR VPWR _705__925/HI _705__925/LO sky130_fd_sc_hd__conb_1
XU$$2212 U$$20/A1 U$$2196/X U$$22/A1 U$$2197/X VGND VGND VPWR VPWR U$$2213/A sky130_fd_sc_hd__a22o_1
XU$$2223 U$$2223/A U$$2257/B VGND VGND VPWR VPWR U$$2223/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_101_2 dadda_fa_4_101_2/A dadda_fa_4_101_2/B dadda_fa_4_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/CIN dadda_fa_5_101_1/CIN sky130_fd_sc_hd__fa_1
XU$$2234 U$$4289/A1 U$$2270/A2 U$$4289/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2235/A
+ sky130_fd_sc_hd__a22o_1
XU$$2245 U$$2245/A U$$2257/B VGND VGND VPWR VPWR U$$2245/X sky130_fd_sc_hd__xor2_1
XFILLER_16_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1500 U$$952/A1 U$$1374/X U$$952/B1 U$$1375/X VGND VGND VPWR VPWR U$$1501/A sky130_fd_sc_hd__a22o_1
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1511 U$$1509/Y _638_/Q _637_/Q U$$1510/X U$$1507/Y VGND VGND VPWR VPWR U$$1511/X
+ sky130_fd_sc_hd__a32o_4
XU$$2256 U$$3900/A1 U$$2270/A2 U$$3489/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2257/A
+ sky130_fd_sc_hd__a22o_1
XU$$2267 U$$2267/A U$$2327/B VGND VGND VPWR VPWR U$$2267/X sky130_fd_sc_hd__xor2_1
XU$$1522 U$$1522/A U$$1614/B VGND VGND VPWR VPWR U$$1522/X sky130_fd_sc_hd__xor2_1
XU$$2278 _591_/Q U$$2326/A2 U$$4335/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2279/A sky130_fd_sc_hd__a22o_1
XFILLER_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1533 U$$26/A1 U$$1591/A2 U$$987/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1534/A sky130_fd_sc_hd__a22o_1
XU$$1544 U$$1544/A U$$1614/B VGND VGND VPWR VPWR U$$1544/X sky130_fd_sc_hd__xor2_1
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2289 U$$2289/A U$$2289/B VGND VGND VPWR VPWR U$$2289/X sky130_fd_sc_hd__xor2_1
XU$$1555 U$$48/A1 U$$1591/A2 U$$50/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1556/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_116_0 _707__927/HI U$$3697/X VGND VGND VPWR VPWR dadda_fa_4_117_2/CIN
+ dadda_ha_3_116_0/SUM sky130_fd_sc_hd__ha_1
XU$$1566 U$$1566/A U$$1580/B VGND VGND VPWR VPWR U$$1566/X sky130_fd_sc_hd__xor2_1
XU$$1577 U$$892/A1 U$$1605/A2 U$$892/B1 U$$1605/B2 VGND VGND VPWR VPWR U$$1578/A sky130_fd_sc_hd__a22o_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1588 U$$1588/A U$$1643/A VGND VGND VPWR VPWR U$$1588/X sky130_fd_sc_hd__xor2_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1599 U$$92/A1 U$$1511/X U$$94/A1 U$$1512/X VGND VGND VPWR VPWR U$$1600/A sky130_fd_sc_hd__a22o_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_115_0 dadda_fa_7_115_0/A dadda_fa_7_115_0/B dadda_fa_7_115_0/CIN VGND
+ VGND VPWR VPWR _540_/D _411_/D sky130_fd_sc_hd__fa_2
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_60_0 dadda_fa_2_60_0/A dadda_fa_2_60_0/B dadda_fa_2_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/B dadda_fa_3_60_2/B sky130_fd_sc_hd__fa_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater400 U$$3977/X VGND VGND VPWR VPWR U$$4045/A2 sky130_fd_sc_hd__buf_12
XFILLER_131_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$207 final_adder.U$$701/A final_adder.U$$573/B1 final_adder.U$$207/B1
+ VGND VGND VPWR VPWR final_adder.U$$207/X sky130_fd_sc_hd__a21o_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater411 U$$3292/X VGND VGND VPWR VPWR U$$3412/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$218 final_adder.U$$713/A final_adder.U$$712/A VGND VGND VPWR VPWR
+ final_adder.U$$300/A sky130_fd_sc_hd__and2_1
Xrepeater422 U$$2607/X VGND VGND VPWR VPWR U$$2729/A2 sky130_fd_sc_hd__buf_12
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$229 final_adder.U$$723/A final_adder.U$$595/B1 final_adder.U$$229/B1
+ VGND VGND VPWR VPWR final_adder.U$$229/X sky130_fd_sc_hd__a21o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater433 U$$2059/X VGND VGND VPWR VPWR U$$2189/A2 sky130_fd_sc_hd__buf_12
Xrepeater444 U$$1511/X VGND VGND VPWR VPWR U$$1591/A2 sky130_fd_sc_hd__buf_12
XFILLER_66_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater455 U$$928/B2 VGND VGND VPWR VPWR U$$910/B2 sky130_fd_sc_hd__buf_12
Xrepeater466 U$$3841/X VGND VGND VPWR VPWR U$$3970/B2 sky130_fd_sc_hd__buf_12
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater477 U$$3156/X VGND VGND VPWR VPWR U$$3253/B2 sky130_fd_sc_hd__buf_12
Xrepeater488 U$$2471/X VGND VGND VPWR VPWR U$$2584/B2 sky130_fd_sc_hd__buf_12
XU$$4170 U$$4170/A1 U$$4114/X U$$4446/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4171/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater499 U$$1923/X VGND VGND VPWR VPWR U$$2052/B2 sky130_fd_sc_hd__buf_12
XU$$4181 U$$4181/A _677_/Q VGND VGND VPWR VPWR U$$4181/X sky130_fd_sc_hd__xor2_1
XU$$4192 U$$630/A1 U$$4114/X U$$632/A1 U$$4115/X VGND VGND VPWR VPWR U$$4193/A sky130_fd_sc_hd__a22o_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3480 U$$3480/A U$$3496/B VGND VGND VPWR VPWR U$$3480/X sky130_fd_sc_hd__xor2_1
XFILLER_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3491 _581_/Q U$$3525/A2 U$$4178/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3492/A sky130_fd_sc_hd__a22o_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2790 U$$50/A1 U$$2796/A2 U$$2790/B1 U$$2826/B2 VGND VGND VPWR VPWR U$$2791/A sky130_fd_sc_hd__a22o_1
XFILLER_22_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_82_1 dadda_fa_4_82_1/A dadda_fa_4_82_1/B dadda_fa_4_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/B dadda_fa_5_82_1/B sky130_fd_sc_hd__fa_1
XFILLER_175_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_75_0 dadda_fa_4_75_0/A dadda_fa_4_75_0/B dadda_fa_4_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/A dadda_fa_5_75_1/A sky130_fd_sc_hd__fa_1
XFILLER_1_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput203 c[51] VGND VGND VPWR VPWR input203/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput214 c[61] VGND VGND VPWR VPWR input214/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput225 c[71] VGND VGND VPWR VPWR input225/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput236 c[81] VGND VGND VPWR VPWR input236/X sky130_fd_sc_hd__clkbuf_1
Xinput247 c[91] VGND VGND VPWR VPWR input247/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$730 final_adder.U$$730/A final_adder.U$$730/B VGND VGND VPWR VPWR
+ _276_/D sky130_fd_sc_hd__xor2_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$741 final_adder.U$$741/A final_adder.U$$741/B VGND VGND VPWR VPWR
+ _287_/D sky130_fd_sc_hd__xor2_1
X_651_ _678_/CLK _651_/D VGND VGND VPWR VPWR _651_/Q sky130_fd_sc_hd__dfxtp_4
XU$$602 U$$54/A1 U$$626/A2 U$$56/A1 U$$553/X VGND VGND VPWR VPWR U$$603/A sky130_fd_sc_hd__a22o_1
XFILLER_56_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$613 U$$613/A U$$661/B VGND VGND VPWR VPWR U$$613/X sky130_fd_sc_hd__xor2_1
XFILLER_29_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$624 U$$76/A1 U$$682/A2 U$$76/B1 U$$553/X VGND VGND VPWR VPWR U$$625/A sky130_fd_sc_hd__a22o_1
X_843__895 VGND VGND VPWR VPWR _843__895/HI U$$819/B1 sky130_fd_sc_hd__conb_1
XU$$635 U$$635/A U$$661/B VGND VGND VPWR VPWR U$$635/X sky130_fd_sc_hd__xor2_1
X_582_ _669_/CLK _582_/D VGND VGND VPWR VPWR _582_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$646 U$$96/B1 U$$682/A2 U$$785/A1 U$$553/X VGND VGND VPWR VPWR U$$647/A sky130_fd_sc_hd__a22o_1
XU$$657 U$$657/A _625_/Q VGND VGND VPWR VPWR U$$657/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$668 U$$942/A1 U$$552/X U$$944/A1 U$$553/X VGND VGND VPWR VPWR U$$669/A sky130_fd_sc_hd__a22o_1
XFILLER_56_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$679 U$$679/A _625_/Q VGND VGND VPWR VPWR U$$679/X sky130_fd_sc_hd__xor2_1
XFILLER_13_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2020 U$$4486/A1 U$$2052/A2 U$$787/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2021/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_32_4 U$$1667/X U$$1800/X U$$1933/X VGND VGND VPWR VPWR dadda_fa_3_33_1/CIN
+ dadda_fa_3_32_3/CIN sky130_fd_sc_hd__fa_1
XU$$2031 U$$2031/A U$$2055/A VGND VGND VPWR VPWR U$$2031/X sky130_fd_sc_hd__xor2_1
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2042 U$$946/A1 U$$2052/A2 U$$948/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2043/A sky130_fd_sc_hd__a22o_1
XFILLER_23_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2053 U$$2053/A U$$2055/A VGND VGND VPWR VPWR U$$2053/X sky130_fd_sc_hd__xor2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2064 U$$2064/A U$$2186/B VGND VGND VPWR VPWR U$$2064/X sky130_fd_sc_hd__xor2_1
XU$$1330 U$$1330/A U$$1336/B VGND VGND VPWR VPWR U$$1330/X sky130_fd_sc_hd__xor2_1
XU$$2075 U$$20/A1 U$$2117/A2 _559_/Q U$$2117/B2 VGND VGND VPWR VPWR U$$2076/A sky130_fd_sc_hd__a22o_1
XU$$1341 U$$930/A1 U$$1341/A2 U$$932/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1342/A sky130_fd_sc_hd__a22o_1
XU$$2086 U$$2086/A U$$2118/B VGND VGND VPWR VPWR U$$2086/X sky130_fd_sc_hd__xor2_1
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2097 U$$3876/B1 U$$2117/A2 U$$4291/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2098/A
+ sky130_fd_sc_hd__a22o_1
XU$$1352 U$$1352/A U$$1369/A VGND VGND VPWR VPWR U$$1352/X sky130_fd_sc_hd__xor2_1
XU$$1363 U$$4514/A1 U$$1367/A2 U$$952/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1364/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1374 U$$1372/Y _636_/Q _635_/Q U$$1373/X U$$1370/Y VGND VGND VPWR VPWR U$$1374/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_188_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1385 U$$1385/A U$$1479/B VGND VGND VPWR VPWR U$$1385/X sky130_fd_sc_hd__xor2_1
XFILLER_148_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1396 U$$26/A1 U$$1474/A2 U$$28/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1397/A sky130_fd_sc_hd__a22o_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_92_0 dadda_fa_5_92_0/A dadda_fa_5_92_0/B dadda_fa_5_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/A dadda_fa_6_92_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_786__838 VGND VGND VPWR VPWR _786__838/HI U$$4417/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_77_6 U$$3752/X U$$3885/X U$$4018/X VGND VGND VPWR VPWR dadda_fa_2_78_2/B
+ dadda_fa_2_77_5/B sky130_fd_sc_hd__fa_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_827__879 VGND VGND VPWR VPWR _827__879/HI U$$4499/B sky130_fd_sc_hd__conb_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$70 _494_/Q _366_/Q VGND VGND VPWR VPWR final_adder.U$$565/B1 final_adder.U$$692/A
+ sky130_fd_sc_hd__ha_1
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$81 _505_/Q _377_/Q VGND VGND VPWR VPWR final_adder.U$$209/B1 final_adder.U$$703/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$92 _516_/Q _388_/Q VGND VGND VPWR VPWR final_adder.U$$587/B1 final_adder.U$$714/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_101_1 input131/X dadda_fa_3_101_1/B dadda_fa_3_101_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_102_0/CIN dadda_fa_4_101_2/A sky130_fd_sc_hd__fa_1
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_122_0 dadda_fa_6_122_0/A dadda_fa_6_122_0/B dadda_fa_6_122_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_123_0/B dadda_fa_7_122_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_103_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_65_4 U$$1733/X U$$1866/X U$$1999/X VGND VGND VPWR VPWR dadda_fa_1_66_6/CIN
+ dadda_fa_1_65_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_42_3 dadda_fa_3_42_3/A dadda_fa_3_42_3/B dadda_fa_3_42_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/B dadda_fa_4_42_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$571 final_adder.U$$698/A final_adder.U$$698/B final_adder.U$$571/B1
+ VGND VGND VPWR VPWR final_adder.U$$699/B sky130_fd_sc_hd__a21o_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_634_ _642_/CLK _634_/D VGND VGND VPWR VPWR _634_/Q sky130_fd_sc_hd__dfxtp_1
XU$$410 _621_/Q VGND VGND VPWR VPWR U$$410/Y sky130_fd_sc_hd__inv_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$421 U$$969/A1 U$$491/A2 U$$971/A1 U$$416/X VGND VGND VPWR VPWR U$$422/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_35_2 dadda_fa_3_35_2/A dadda_fa_3_35_2/B dadda_fa_3_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/A dadda_fa_4_35_2/B sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$593 final_adder.U$$720/A final_adder.U$$720/B final_adder.U$$593/B1
+ VGND VGND VPWR VPWR final_adder.U$$721/B sky130_fd_sc_hd__a21o_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$432 U$$432/A U$$530/B VGND VGND VPWR VPWR U$$432/X sky130_fd_sc_hd__xor2_1
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$443 U$$32/A1 U$$545/A2 U$$34/A1 U$$416/X VGND VGND VPWR VPWR U$$444/A sky130_fd_sc_hd__a22o_1
XFILLER_45_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$454 U$$454/A U$$530/B VGND VGND VPWR VPWR U$$454/X sky130_fd_sc_hd__xor2_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_1 U$$1925/X U$$2021/B input177/X VGND VGND VPWR VPWR dadda_fa_4_29_0/CIN
+ dadda_fa_4_28_2/A sky130_fd_sc_hd__fa_2
XU$$465 U$$54/A1 U$$545/A2 U$$56/A1 U$$416/X VGND VGND VPWR VPWR U$$466/A sky130_fd_sc_hd__a22o_1
X_565_ _576_/CLK _565_/D VGND VGND VPWR VPWR _565_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$476 U$$476/A U$$547/A VGND VGND VPWR VPWR U$$476/X sky130_fd_sc_hd__xor2_1
XU$$487 U$$759/B1 U$$491/A2 U$$78/A1 U$$416/X VGND VGND VPWR VPWR U$$488/A sky130_fd_sc_hd__a22o_1
XFILLER_60_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$498 U$$498/A U$$547/A VGND VGND VPWR VPWR U$$498/X sky130_fd_sc_hd__xor2_1
X_496_ _496_/CLK _496_/D VGND VGND VPWR VPWR _496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_87_5 dadda_fa_2_87_5/A dadda_fa_2_87_5/B dadda_fa_2_87_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_2/A dadda_fa_4_87_0/A sky130_fd_sc_hd__fa_2
XFILLER_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_30_1 U$$466/X U$$599/X U$$732/X VGND VGND VPWR VPWR dadda_fa_3_31_1/B
+ dadda_fa_3_30_3/A sky130_fd_sc_hd__fa_1
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1160 U$$64/A1 U$$1200/A2 U$$66/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1161/A sky130_fd_sc_hd__a22o_1
XFILLER_149_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1171 U$$1171/A U$$1189/B VGND VGND VPWR VPWR U$$1171/X sky130_fd_sc_hd__xor2_1
XFILLER_189_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1182 U$$908/A1 U$$1218/A2 U$$88/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1183/A sky130_fd_sc_hd__a22o_1
XU$$1193 U$$1193/A U$$1232/A VGND VGND VPWR VPWR U$$1193/X sky130_fd_sc_hd__xor2_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_117_1 dadda_fa_5_117_1/A dadda_fa_5_117_1/B dadda_fa_5_117_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/B dadda_fa_7_117_0/A sky130_fd_sc_hd__fa_2
XFILLER_176_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_82_4 U$$2831/X U$$2964/X U$$3097/X VGND VGND VPWR VPWR dadda_fa_2_83_2/CIN
+ dadda_fa_2_82_5/A sky130_fd_sc_hd__fa_2
XFILLER_160_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_75_3 U$$2817/X U$$2950/X U$$3083/X VGND VGND VPWR VPWR dadda_fa_2_76_1/B
+ dadda_fa_2_75_4/B sky130_fd_sc_hd__fa_1
XFILLER_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_52_2 dadda_fa_4_52_2/A dadda_fa_4_52_2/B dadda_fa_4_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/CIN dadda_fa_5_52_1/CIN sky130_fd_sc_hd__fa_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_2 U$$3335/X U$$3468/X U$$3601/X VGND VGND VPWR VPWR dadda_fa_2_69_1/A
+ dadda_fa_2_68_4/A sky130_fd_sc_hd__fa_2
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_45_1 dadda_fa_4_45_1/A dadda_fa_4_45_1/B dadda_fa_4_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/B dadda_fa_5_45_1/B sky130_fd_sc_hd__fa_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_22_0 dadda_fa_7_22_0/A dadda_fa_7_22_0/B dadda_fa_7_22_0/CIN VGND VGND
+ VPWR VPWR _447_/D _318_/D sky130_fd_sc_hd__fa_2
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_0 dadda_fa_4_38_0/A dadda_fa_4_38_0/B dadda_fa_4_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/A dadda_fa_5_38_1/A sky130_fd_sc_hd__fa_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _483_/CLK _350_/D VGND VGND VPWR VPWR _350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_281_ _612_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_0_57_2 U$$919/X U$$1052/X VGND VGND VPWR VPWR dadda_fa_1_58_7/CIN dadda_fa_2_57_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_190_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_70_2 U$$1211/X U$$1344/X U$$1477/X VGND VGND VPWR VPWR dadda_fa_1_71_7/A
+ dadda_fa_1_70_8/B sky130_fd_sc_hd__fa_1
XFILLER_118_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_63_1 U$$532/X U$$665/X U$$798/X VGND VGND VPWR VPWR dadda_fa_1_64_5/CIN
+ dadda_fa_1_63_7/CIN sky130_fd_sc_hd__fa_2
XFILLER_49_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_40_0 dadda_fa_3_40_0/A dadda_fa_3_40_0/B dadda_fa_3_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/B dadda_fa_4_40_1/CIN sky130_fd_sc_hd__fa_2
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_0 U$$119/X U$$252/X U$$385/X VGND VGND VPWR VPWR dadda_fa_1_57_7/B
+ dadda_fa_1_56_8/B sky130_fd_sc_hd__fa_2
XFILLER_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$240 U$$240/A U$$274/A VGND VGND VPWR VPWR U$$240/X sky130_fd_sc_hd__xor2_1
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_617_ _621_/CLK _617_/D VGND VGND VPWR VPWR _617_/Q sky130_fd_sc_hd__dfxtp_4
XU$$251 U$$799/A1 U$$141/X U$$938/A1 U$$142/X VGND VGND VPWR VPWR U$$252/A sky130_fd_sc_hd__a22o_1
XFILLER_45_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$262 U$$262/A U$$262/B VGND VGND VPWR VPWR U$$262/X sky130_fd_sc_hd__xor2_2
XU$$273 _619_/Q VGND VGND VPWR VPWR U$$273/Y sky130_fd_sc_hd__inv_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$284 U$$8/B1 U$$278/X U$$12/A1 U$$279/X VGND VGND VPWR VPWR U$$285/A sky130_fd_sc_hd__a22o_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$295 U$$295/A U$$391/B VGND VGND VPWR VPWR U$$295/X sky130_fd_sc_hd__xor2_1
X_548_ _656_/CLK _548_/D VGND VGND VPWR VPWR _548_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_479_ _480_/CLK _479_/D VGND VGND VPWR VPWR _479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1 U$$1/A VGND VGND VPWR VPWR U$$3/B sky130_fd_sc_hd__inv_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$9 _433_/Q _305_/Q VGND VGND VPWR VPWR final_adder.U$$9/COUT final_adder.U$$9/SUM
+ sky130_fd_sc_hd__ha_2
Xoutput304 _195_/Q VGND VGND VPWR VPWR o[27] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_3 U$$4181/X U$$4314/X U$$4447/X VGND VGND VPWR VPWR dadda_fa_3_93_1/B
+ dadda_fa_3_92_3/B sky130_fd_sc_hd__fa_1
Xoutput315 _205_/Q VGND VGND VPWR VPWR o[37] sky130_fd_sc_hd__buf_2
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput326 _215_/Q VGND VGND VPWR VPWR o[47] sky130_fd_sc_hd__buf_2
XFILLER_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput337 _225_/Q VGND VGND VPWR VPWR o[57] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_2 dadda_fa_2_85_2/A dadda_fa_2_85_2/B dadda_fa_2_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/A dadda_fa_3_85_3/A sky130_fd_sc_hd__fa_2
Xoutput348 _235_/Q VGND VGND VPWR VPWR o[67] sky130_fd_sc_hd__buf_2
Xoutput359 _245_/Q VGND VGND VPWR VPWR o[77] sky130_fd_sc_hd__buf_2
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_62_1 dadda_fa_5_62_1/A dadda_fa_5_62_1/B dadda_fa_5_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/B dadda_fa_7_62_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_78_1 dadda_fa_2_78_1/A dadda_fa_2_78_1/B dadda_fa_2_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/CIN dadda_fa_3_78_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_55_0 dadda_fa_5_55_0/A dadda_fa_5_55_0/B dadda_fa_5_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/A dadda_fa_6_55_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_84_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_8 input206/X dadda_fa_1_54_8/B dadda_fa_1_54_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_55_3/A dadda_fa_3_54_0/A sky130_fd_sc_hd__fa_2
XFILLER_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_101_0 U$$2602/Y U$$2736/X U$$2869/X VGND VGND VPWR VPWR dadda_fa_3_102_1/CIN
+ dadda_fa_3_101_3/A sky130_fd_sc_hd__fa_1
XFILLER_51_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_80_1 U$$1497/X U$$1630/X U$$1763/X VGND VGND VPWR VPWR dadda_fa_2_81_1/A
+ dadda_fa_2_80_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_133_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_0 U$$1882/X U$$2015/X U$$2148/X VGND VGND VPWR VPWR dadda_fa_2_74_0/B
+ dadda_fa_2_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_150_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3309 U$$3309/A U$$3413/B VGND VGND VPWR VPWR U$$3309/X sky130_fd_sc_hd__xor2_1
XFILLER_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2608 U$$2606/B U$$2603/A _654_/Q U$$2603/Y VGND VGND VPWR VPWR U$$2608/X sky130_fd_sc_hd__a22o_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2619 U$$14/B1 U$$2667/A2 U$$4265/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2620/A sky130_fd_sc_hd__a22o_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1907 U$$948/A1 U$$1785/X U$$950/A1 U$$1786/X VGND VGND VPWR VPWR U$$1908/A sky130_fd_sc_hd__a22o_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1918 U$$1918/A VGND VGND VPWR VPWR U$$1918/Y sky130_fd_sc_hd__inv_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _543_/CLK _402_/D VGND VGND VPWR VPWR _402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1929 U$$1929/A U$$2021/B VGND VGND VPWR VPWR U$$1929/X sky130_fd_sc_hd__xor2_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_333_ _333_/CLK _333_/D VGND VGND VPWR VPWR _333_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_264_ _280_/CLK _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ _329_/CLK _195_/D VGND VGND VPWR VPWR _195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_95_1 dadda_fa_3_95_1/A dadda_fa_3_95_1/B dadda_fa_3_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/CIN dadda_fa_4_95_2/A sky130_fd_sc_hd__fa_2
XFILLER_115_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_72_0 dadda_fa_6_72_0/A dadda_fa_6_72_0/B dadda_fa_6_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_73_0/B dadda_fa_7_72_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_88_0 dadda_fa_3_88_0/A dadda_fa_3_88_0/B dadda_fa_3_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/B dadda_fa_4_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4500 U$$4500/A1 U$$4388/X U$$4502/A1 U$$4389/X VGND VGND VPWR VPWR U$$4501/A sky130_fd_sc_hd__a22o_1
XU$$4511 U$$4511/A U$$4511/B VGND VGND VPWR VPWR U$$4511/X sky130_fd_sc_hd__xor2_2
XFILLER_110_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$14 U$$14/A1 U$$4/X U$$14/B1 U$$5/X VGND VGND VPWR VPWR U$$15/A sky130_fd_sc_hd__a22o_1
XU$$25 U$$25/A U$$89/B VGND VGND VPWR VPWR U$$25/X sky130_fd_sc_hd__xor2_1
XU$$3810 U$$3810/A U$$3835/A VGND VGND VPWR VPWR U$$3810/X sky130_fd_sc_hd__xor2_1
XU$$3821 U$$4506/A1 U$$3703/X U$$4508/A1 U$$3704/X VGND VGND VPWR VPWR U$$3822/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_117_0 U$$3698/Y U$$3832/X U$$3965/X VGND VGND VPWR VPWR dadda_fa_5_118_0/A
+ dadda_fa_5_117_1/A sky130_fd_sc_hd__fa_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$36 U$$36/A1 U$$4/X U$$38/A1 U$$5/X VGND VGND VPWR VPWR U$$37/A sky130_fd_sc_hd__a22o_1
XU$$3832 U$$3832/A U$$3835/A VGND VGND VPWR VPWR U$$3832/X sky130_fd_sc_hd__xor2_1
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$47 U$$47/A U$$3/A VGND VGND VPWR VPWR U$$47/X sky130_fd_sc_hd__xor2_1
XFILLER_65_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3843 U$$3843/A U$$3893/B VGND VGND VPWR VPWR U$$3843/X sky130_fd_sc_hd__xor2_1
XU$$58 U$$58/A1 U$$4/X U$$60/A1 U$$5/X VGND VGND VPWR VPWR U$$59/A sky130_fd_sc_hd__a22o_1
XU$$69 U$$69/A U$$9/B VGND VGND VPWR VPWR U$$69/X sky130_fd_sc_hd__xor2_1
XU$$3854 U$$975/B1 U$$3840/X U$$979/A1 U$$3841/X VGND VGND VPWR VPWR U$$3855/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_5_4_0 U$$15/X U$$148/X VGND VGND VPWR VPWR dadda_fa_6_5_0/CIN dadda_fa_7_4_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_92_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3865 U$$3865/A U$$3893/B VGND VGND VPWR VPWR U$$3865/X sky130_fd_sc_hd__xor2_1
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3876 U$$4424/A1 U$$3912/A2 U$$3876/B1 U$$3912/B2 VGND VGND VPWR VPWR U$$3877/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3887 U$$3887/A U$$3929/B VGND VGND VPWR VPWR U$$3887/X sky130_fd_sc_hd__xor2_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3898 U$$4446/A1 U$$3970/A2 _580_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3899/A sky130_fd_sc_hd__a22o_1
XFILLER_36_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_90_0 U$$3246/X U$$3379/X U$$3512/X VGND VGND VPWR VPWR dadda_fa_3_91_0/B
+ dadda_fa_3_90_2/B sky130_fd_sc_hd__fa_2
XFILLER_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_46_6 U$$2493/X U$$2626/X VGND VGND VPWR VPWR dadda_fa_2_47_3/CIN dadda_fa_3_46_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_5 U$$2372/X U$$2505/X U$$2638/X VGND VGND VPWR VPWR dadda_fa_2_53_2/A
+ dadda_fa_2_52_5/A sky130_fd_sc_hd__fa_2
XFILLER_110_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_45_4 U$$1693/X U$$1826/X U$$1959/X VGND VGND VPWR VPWR dadda_fa_2_46_3/B
+ dadda_fa_2_45_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_83_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_15_2 input163/X dadda_fa_4_15_2/B dadda_ha_3_15_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_5_16_0/CIN dadda_fa_5_15_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_52_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3106 U$$4476/A1 U$$3146/A2 U$$94/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3107/A sky130_fd_sc_hd__a22o_1
XFILLER_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3117 U$$3117/A U$$3137/B VGND VGND VPWR VPWR U$$3117/X sky130_fd_sc_hd__xor2_1
XFILLER_143_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3128 _605_/Q U$$3018/X _606_/Q U$$3019/X VGND VGND VPWR VPWR U$$3129/A sky130_fd_sc_hd__a22o_1
XU$$3139 U$$3139/A _661_/Q VGND VGND VPWR VPWR U$$3139/X sky130_fd_sc_hd__xor2_1
XU$$2405 U$$2953/A1 U$$2421/A2 U$$76/B1 U$$2421/B2 VGND VGND VPWR VPWR U$$2406/A sky130_fd_sc_hd__a22o_1
XU$$2416 U$$2416/A U$$2436/B VGND VGND VPWR VPWR U$$2416/X sky130_fd_sc_hd__xor2_1
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2427 U$$98/A1 U$$2463/A2 U$$98/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2428/A sky130_fd_sc_hd__a22o_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2438 U$$2438/A U$$2464/B VGND VGND VPWR VPWR U$$2438/X sky130_fd_sc_hd__xor2_1
XU$$1704 U$$60/A1 U$$1726/A2 U$$4446/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1705/A sky130_fd_sc_hd__a22o_1
XU$$2449 U$$942/A1 U$$2463/A2 U$$4506/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2450/A
+ sky130_fd_sc_hd__a22o_1
XU$$1715 U$$1715/A U$$1739/B VGND VGND VPWR VPWR U$$1715/X sky130_fd_sc_hd__xor2_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1726 U$$902/B1 U$$1726/A2 U$$84/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1727/A sky130_fd_sc_hd__a22o_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1737 U$$1737/A _641_/Q VGND VGND VPWR VPWR U$$1737/X sky130_fd_sc_hd__xor2_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1748 U$$926/A1 U$$1770/A2 U$$928/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1749/A sky130_fd_sc_hd__a22o_1
XFILLER_159_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1759 U$$1759/A _641_/Q VGND VGND VPWR VPWR U$$1759/X sky130_fd_sc_hd__xor2_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_316_ _461_/CLK _316_/D VGND VGND VPWR VPWR _316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ _501_/CLK _247_/D VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_1
Xinput14 a[21] VGND VGND VPWR VPWR _637_/D sky130_fd_sc_hd__buf_2
Xinput25 a[31] VGND VGND VPWR VPWR _647_/D sky130_fd_sc_hd__clkbuf_4
Xinput36 a[41] VGND VGND VPWR VPWR _657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput47 a[51] VGND VGND VPWR VPWR _667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput58 a[61] VGND VGND VPWR VPWR _677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_178_ _464_/CLK _178_/D VGND VGND VPWR VPWR _178_/Q sky130_fd_sc_hd__dfxtp_2
Xinput69 b[13] VGND VGND VPWR VPWR _565_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_182_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_62_4 dadda_fa_2_62_4/A dadda_fa_2_62_4/B dadda_fa_2_62_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/CIN dadda_fa_3_62_3/CIN sky130_fd_sc_hd__fa_2
Xrepeater604 U$$391/B VGND VGND VPWR VPWR U$$357/B sky130_fd_sc_hd__buf_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater615 _614_/Q VGND VGND VPWR VPWR U$$4379/A1 sky130_fd_sc_hd__buf_12
Xrepeater626 U$$4504/A1 VGND VGND VPWR VPWR U$$942/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater637 _603_/Q VGND VGND VPWR VPWR U$$4494/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_55_3 dadda_fa_2_55_3/A dadda_fa_2_55_3/B dadda_fa_2_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/B dadda_fa_3_55_3/B sky130_fd_sc_hd__fa_2
Xrepeater648 _598_/Q VGND VGND VPWR VPWR U$$785/A1 sky130_fd_sc_hd__buf_12
XU$$4330 U$$4330/A U$$4384/A VGND VGND VPWR VPWR U$$4330/X sky130_fd_sc_hd__xor2_1
XU$$4341 U$$94/A1 U$$4377/A2 U$$94/B1 U$$4377/B2 VGND VGND VPWR VPWR U$$4342/A sky130_fd_sc_hd__a22o_1
Xrepeater659 _593_/Q VGND VGND VPWR VPWR U$$90/A1 sky130_fd_sc_hd__buf_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4352 U$$4352/A U$$4384/A VGND VGND VPWR VPWR U$$4352/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_2 dadda_fa_2_48_2/A dadda_fa_2_48_2/B dadda_fa_2_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/A dadda_fa_3_48_3/A sky130_fd_sc_hd__fa_1
XU$$4363 U$$4500/A1 U$$4377/A2 U$$4502/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4364/A
+ sky130_fd_sc_hd__a22o_1
XU$$4374 U$$4374/A U$$4384/A VGND VGND VPWR VPWR U$$4374/X sky130_fd_sc_hd__xor2_1
XU$$3640 _587_/Q U$$3668/A2 _588_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3641/A sky130_fd_sc_hd__a22o_1
XU$$4385 U$$4385/A VGND VGND VPWR VPWR U$$4387/B sky130_fd_sc_hd__inv_1
XFILLER_77_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4396 _554_/Q U$$4388/X _555_/Q U$$4389/X VGND VGND VPWR VPWR U$$4397/A sky130_fd_sc_hd__a22o_1
XU$$3651 U$$3651/A U$$3698/A VGND VGND VPWR VPWR U$$3651/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_25_1 dadda_fa_5_25_1/A dadda_fa_5_25_1/B dadda_fa_5_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/B dadda_fa_7_25_0/A sky130_fd_sc_hd__fa_1
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3662 U$$4484/A1 U$$3668/A2 _599_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3663/A sky130_fd_sc_hd__a22o_1
XU$$3673 U$$3673/A _669_/Q VGND VGND VPWR VPWR U$$3673/X sky130_fd_sc_hd__xor2_1
XU$$3684 U$$4506/A1 U$$3566/X U$$4508/A1 U$$3567/X VGND VGND VPWR VPWR U$$3685/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_18_0 dadda_fa_5_18_0/A dadda_fa_5_18_0/B dadda_fa_5_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/A dadda_fa_6_18_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_46_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2950 U$$2950/A U$$2960/B VGND VGND VPWR VPWR U$$2950/X sky130_fd_sc_hd__xor2_1
XU$$3695 U$$3695/A U$$3698/A VGND VGND VPWR VPWR U$$3695/X sky130_fd_sc_hd__xor2_1
XFILLER_34_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2961 _590_/Q U$$2975/A2 U$$908/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2962/A sky130_fd_sc_hd__a22o_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2972 U$$2972/A _659_/Q VGND VGND VPWR VPWR U$$2972/X sky130_fd_sc_hd__xor2_1
XU$$2983 _601_/Q U$$2881/X _602_/Q U$$2882/X VGND VGND VPWR VPWR U$$2984/A sky130_fd_sc_hd__a22o_1
XFILLER_61_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2994 U$$2994/A U$$2996/B VGND VGND VPWR VPWR U$$2994/X sky130_fd_sc_hd__xor2_1
XFILLER_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_50_2 U$$905/X U$$1038/X U$$1171/X VGND VGND VPWR VPWR dadda_fa_2_51_1/A
+ dadda_fa_2_50_4/A sky130_fd_sc_hd__fa_1
XFILLER_21_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$806 U$$806/A U$$822/A VGND VGND VPWR VPWR U$$806/X sky130_fd_sc_hd__xor2_1
XU$$817 U$$952/B1 U$$817/A2 U$$956/A1 U$$817/B2 VGND VGND VPWR VPWR U$$818/A sky130_fd_sc_hd__a22o_1
XFILLER_113_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_43_1 U$$492/X U$$625/X U$$758/X VGND VGND VPWR VPWR dadda_fa_2_44_3/A
+ dadda_fa_2_43_5/A sky130_fd_sc_hd__fa_1
XU$$828 U$$828/A1 U$$910/A2 U$$8/A1 U$$910/B2 VGND VGND VPWR VPWR U$$829/A sky130_fd_sc_hd__a22o_1
XU$$839 U$$839/A U$$959/A VGND VGND VPWR VPWR U$$839/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_20_0 U$$1479/B input169/X dadda_fa_4_20_0/CIN VGND VGND VPWR VPWR dadda_fa_5_21_0/A
+ dadda_fa_5_20_1/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_36_0 U$$79/X U$$212/X U$$345/X VGND VGND VPWR VPWR dadda_fa_2_37_5/A dadda_fa_2_36_5/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_189_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_72_3 dadda_fa_3_72_3/A dadda_fa_3_72_3/B dadda_fa_3_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/B dadda_fa_4_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_65_2 dadda_fa_3_65_2/A dadda_fa_3_65_2/B dadda_fa_3_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/A dadda_fa_4_65_2/B sky130_fd_sc_hd__fa_1
XFILLER_117_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_58_1 dadda_fa_3_58_1/A dadda_fa_3_58_1/B dadda_fa_3_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/CIN dadda_fa_4_58_2/A sky130_fd_sc_hd__fa_1
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_35_0 dadda_fa_6_35_0/A dadda_fa_6_35_0/B dadda_fa_6_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_36_0/B dadda_fa_7_35_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2202 _553_/Q U$$2270/A2 U$$4122/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2203/A sky130_fd_sc_hd__a22o_1
XU$$2213 U$$2213/A U$$2289/B VGND VGND VPWR VPWR U$$2213/X sky130_fd_sc_hd__xor2_1
XU$$2224 U$$30/B1 U$$2270/A2 U$$3457/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2225/A sky130_fd_sc_hd__a22o_1
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2235 U$$2235/A U$$2257/B VGND VGND VPWR VPWR U$$2235/X sky130_fd_sc_hd__xor2_1
XU$$1501 U$$1501/A _637_/Q VGND VGND VPWR VPWR U$$1501/X sky130_fd_sc_hd__xor2_1
XU$$2246 U$$876/A1 U$$2270/A2 U$$878/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2247/A sky130_fd_sc_hd__a22o_1
XU$$1512 U$$1510/B _637_/Q _638_/Q U$$1507/Y VGND VGND VPWR VPWR U$$1512/X sky130_fd_sc_hd__a22o_4
XFILLER_90_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2257 U$$2257/A U$$2257/B VGND VGND VPWR VPWR U$$2257/X sky130_fd_sc_hd__xor2_1
XU$$2268 U$$759/B1 U$$2196/X U$$78/A1 U$$2197/X VGND VGND VPWR VPWR U$$2269/A sky130_fd_sc_hd__a22o_1
XU$$1523 U$$14/B1 U$$1591/A2 U$$18/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1524/A sky130_fd_sc_hd__a22o_1
XU$$2279 U$$2279/A U$$2289/B VGND VGND VPWR VPWR U$$2279/X sky130_fd_sc_hd__xor2_1
XU$$1534 U$$1534/A U$$1580/B VGND VGND VPWR VPWR U$$1534/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1545 U$$38/A1 U$$1591/A2 U$$3191/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1546/A sky130_fd_sc_hd__a22o_1
XU$$1556 U$$1556/A U$$1580/B VGND VGND VPWR VPWR U$$1556/X sky130_fd_sc_hd__xor2_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1567 _578_/Q U$$1591/A2 U$$4446/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1568/A sky130_fd_sc_hd__a22o_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1578 U$$1578/A U$$1580/B VGND VGND VPWR VPWR U$$1578/X sky130_fd_sc_hd__xor2_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1589 U$$630/A1 U$$1591/A2 U$$84/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1590/A sky130_fd_sc_hd__a22o_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_108_0 dadda_fa_7_108_0/A dadda_fa_7_108_0/B dadda_fa_7_108_0/CIN VGND
+ VGND VPWR VPWR _533_/D _404_/D sky130_fd_sc_hd__fa_2
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_1 dadda_fa_2_60_1/A dadda_fa_2_60_1/B dadda_fa_2_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/CIN dadda_fa_3_60_2/CIN sky130_fd_sc_hd__fa_2
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater401 U$$3840/X VGND VGND VPWR VPWR U$$3912/A2 sky130_fd_sc_hd__buf_12
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$208 final_adder.U$$703/A final_adder.U$$702/A VGND VGND VPWR VPWR
+ final_adder.U$$296/B sky130_fd_sc_hd__and2_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater412 U$$3155/X VGND VGND VPWR VPWR U$$3243/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$219 final_adder.U$$713/A final_adder.U$$585/B1 final_adder.U$$219/B1
+ VGND VGND VPWR VPWR final_adder.U$$219/X sky130_fd_sc_hd__a21o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater423 U$$2574/A2 VGND VGND VPWR VPWR U$$2534/A2 sky130_fd_sc_hd__buf_12
Xrepeater434 U$$2048/A2 VGND VGND VPWR VPWR U$$2036/A2 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_53_0 dadda_fa_2_53_0/A dadda_fa_2_53_0/B dadda_fa_2_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/B dadda_fa_3_53_2/B sky130_fd_sc_hd__fa_2
Xrepeater445 U$$1511/X VGND VGND VPWR VPWR U$$1641/A2 sky130_fd_sc_hd__buf_12
XFILLER_111_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater456 U$$827/X VGND VGND VPWR VPWR U$$928/B2 sky130_fd_sc_hd__buf_12
Xrepeater467 U$$3704/X VGND VGND VPWR VPWR U$$3783/B2 sky130_fd_sc_hd__buf_12
Xrepeater478 U$$3146/B2 VGND VGND VPWR VPWR U$$3090/B2 sky130_fd_sc_hd__buf_12
XU$$4160 _573_/Q U$$4198/A2 _574_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4161/A sky130_fd_sc_hd__a22o_1
XFILLER_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater489 U$$2463/B2 VGND VGND VPWR VPWR U$$2421/B2 sky130_fd_sc_hd__buf_12
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4171 U$$4171/A U$$4197/B VGND VGND VPWR VPWR U$$4171/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4182 U$$70/B1 U$$4244/A2 U$$759/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4183/A sky130_fd_sc_hd__a22o_1
XU$$4193 U$$4193/A U$$4247/A VGND VGND VPWR VPWR U$$4193/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3470 U$$3470/A U$$3496/B VGND VGND VPWR VPWR U$$3470/X sky130_fd_sc_hd__xor2_1
XU$$3481 U$$4303/A1 U$$3525/A2 U$$4442/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3482/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3492 U$$3492/A U$$3496/B VGND VGND VPWR VPWR U$$3492/X sky130_fd_sc_hd__xor2_1
XFILLER_53_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2780 U$$4424/A1 U$$2796/A2 U$$4289/A1 U$$2834/B2 VGND VGND VPWR VPWR U$$2781/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_7_0 U$$21/X U$$154/X U$$287/X VGND VGND VPWR VPWR dadda_fa_6_8_0/A dadda_fa_6_7_0/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2791 U$$2791/A U$$2797/B VGND VGND VPWR VPWR U$$2791/X sky130_fd_sc_hd__xor2_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_82_2 dadda_fa_4_82_2/A dadda_fa_4_82_2/B dadda_fa_4_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/CIN dadda_fa_5_82_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_75_1 dadda_fa_4_75_1/A dadda_fa_4_75_1/B dadda_fa_4_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/B dadda_fa_5_75_1/B sky130_fd_sc_hd__fa_1
XFILLER_136_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_687__907 VGND VGND VPWR VPWR _687__907/HI _687__907/LO sky130_fd_sc_hd__conb_1
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_52_0 dadda_fa_7_52_0/A dadda_fa_7_52_0/B dadda_fa_7_52_0/CIN VGND VGND
+ VPWR VPWR _477_/D _348_/D sky130_fd_sc_hd__fa_2
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_68_0 dadda_fa_4_68_0/A dadda_fa_4_68_0/B dadda_fa_4_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/A dadda_fa_5_68_1/A sky130_fd_sc_hd__fa_1
Xinput204 c[52] VGND VGND VPWR VPWR input204/X sky130_fd_sc_hd__buf_2
XFILLER_0_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput215 c[62] VGND VGND VPWR VPWR input215/X sky130_fd_sc_hd__buf_2
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput226 c[72] VGND VGND VPWR VPWR input226/X sky130_fd_sc_hd__buf_2
Xinput237 c[82] VGND VGND VPWR VPWR input237/X sky130_fd_sc_hd__clkbuf_2
Xinput248 c[92] VGND VGND VPWR VPWR input248/X sky130_fd_sc_hd__buf_2
Xfinal_adder.U$$720 final_adder.U$$720/A final_adder.U$$720/B VGND VGND VPWR VPWR
+ _266_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$731 final_adder.U$$731/A final_adder.U$$731/B VGND VGND VPWR VPWR
+ _277_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$742 final_adder.U$$742/A final_adder.U$$742/B VGND VGND VPWR VPWR
+ _288_/D sky130_fd_sc_hd__xor2_2
XFILLER_29_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_650_ _650_/CLK _650_/D VGND VGND VPWR VPWR _650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$603 U$$603/A U$$623/B VGND VGND VPWR VPWR U$$603/X sky130_fd_sc_hd__xor2_1
XFILLER_112_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$614 U$$66/A1 U$$626/A2 U$$68/A1 U$$553/X VGND VGND VPWR VPWR U$$615/A sky130_fd_sc_hd__a22o_1
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$625 U$$625/A U$$661/B VGND VGND VPWR VPWR U$$625/X sky130_fd_sc_hd__xor2_1
XFILLER_84_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$636 U$$88/A1 U$$682/A2 U$$90/A1 U$$553/X VGND VGND VPWR VPWR U$$637/A sky130_fd_sc_hd__a22o_1
X_581_ _581_/CLK _581_/D VGND VGND VPWR VPWR _581_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$647 U$$647/A U$$661/B VGND VGND VPWR VPWR U$$647/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$658 _603_/Q U$$682/A2 U$$934/A1 U$$553/X VGND VGND VPWR VPWR U$$659/A sky130_fd_sc_hd__a22o_1
XU$$669 U$$669/A _625_/Q VGND VGND VPWR VPWR U$$669/X sky130_fd_sc_hd__xor2_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_70_0 dadda_fa_3_70_0/A dadda_fa_3_70_0/B dadda_fa_3_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/B dadda_fa_4_70_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2010 U$$914/A1 U$$2036/A2 U$$92/B1 U$$2036/B2 VGND VGND VPWR VPWR U$$2011/A sky130_fd_sc_hd__a22o_1
XU$$2021 U$$2021/A U$$2021/B VGND VGND VPWR VPWR U$$2021/X sky130_fd_sc_hd__xor2_1
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2032 U$$799/A1 U$$2048/A2 U$$938/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$2033/A sky130_fd_sc_hd__a22o_1
XU$$2043 U$$2043/A U$$2055/A VGND VGND VPWR VPWR U$$2043/X sky130_fd_sc_hd__xor2_1
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2054 U$$2055/A VGND VGND VPWR VPWR U$$2054/Y sky130_fd_sc_hd__inv_1
XU$$2065 U$$8/B1 U$$2117/A2 U$$971/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2066/A sky130_fd_sc_hd__a22o_1
XU$$1320 U$$1320/A U$$1369/A VGND VGND VPWR VPWR U$$1320/X sky130_fd_sc_hd__xor2_1
XU$$1331 U$$98/A1 U$$1237/X U$$98/B1 U$$1238/X VGND VGND VPWR VPWR U$$1332/A sky130_fd_sc_hd__a22o_1
XFILLER_90_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2076 U$$2076/A U$$2186/B VGND VGND VPWR VPWR U$$2076/X sky130_fd_sc_hd__xor2_1
XU$$2087 U$$30/B1 U$$2117/A2 U$$3457/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2088/A sky130_fd_sc_hd__a22o_1
XU$$1342 U$$1342/A U$$1342/B VGND VGND VPWR VPWR U$$1342/X sky130_fd_sc_hd__xor2_1
XFILLER_90_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2098 U$$2098/A U$$2118/B VGND VGND VPWR VPWR U$$2098/X sky130_fd_sc_hd__xor2_1
XU$$1353 _608_/Q U$$1367/A2 _609_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1354/A sky130_fd_sc_hd__a22o_1
XU$$1364 U$$1364/A _635_/Q VGND VGND VPWR VPWR U$$1364/X sky130_fd_sc_hd__xor2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1375 U$$1373/B _635_/Q _636_/Q U$$1370/Y VGND VGND VPWR VPWR U$$1375/X sky130_fd_sc_hd__a22o_4
XFILLER_43_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1386 U$$14/B1 U$$1474/A2 U$$18/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1387/A sky130_fd_sc_hd__a22o_1
XFILLER_31_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1397 U$$1397/A U$$1479/B VGND VGND VPWR VPWR U$$1397/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_92_1 dadda_fa_5_92_1/A dadda_fa_5_92_1/B dadda_fa_5_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/B dadda_fa_7_92_0/A sky130_fd_sc_hd__fa_1
XFILLER_11_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_85_0 dadda_fa_5_85_0/A dadda_fa_5_85_0/B dadda_fa_5_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/A dadda_fa_6_85_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_77_7 U$$4151/X U$$4284/X U$$4417/X VGND VGND VPWR VPWR dadda_fa_2_78_2/CIN
+ dadda_fa_2_77_5/CIN sky130_fd_sc_hd__fa_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$60 _484_/Q _356_/Q VGND VGND VPWR VPWR final_adder.U$$555/B1 final_adder.U$$682/A
+ sky130_fd_sc_hd__ha_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$71 _495_/Q _367_/Q VGND VGND VPWR VPWR final_adder.U$$199/B1 final_adder.U$$693/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$82 _506_/Q _378_/Q VGND VGND VPWR VPWR final_adder.U$$577/B1 final_adder.U$$704/A
+ sky130_fd_sc_hd__ha_1
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$93 _517_/Q _389_/Q VGND VGND VPWR VPWR final_adder.U$$221/B1 final_adder.U$$715/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_101_2 dadda_fa_3_101_2/A dadda_fa_3_101_2/B dadda_fa_3_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/A dadda_fa_4_101_2/B sky130_fd_sc_hd__fa_1
XFILLER_163_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_810__862 VGND VGND VPWR VPWR _810__862/HI U$$4465/B sky130_fd_sc_hd__conb_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_65_5 U$$2132/X U$$2265/X U$$2398/X VGND VGND VPWR VPWR dadda_fa_1_66_7/A
+ dadda_fa_2_65_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_6_115_0 dadda_fa_6_115_0/A dadda_fa_6_115_0/B dadda_fa_6_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_116_0/B dadda_fa_7_115_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$561 final_adder.U$$688/A final_adder.U$$688/B final_adder.U$$561/B1
+ VGND VGND VPWR VPWR final_adder.U$$689/B sky130_fd_sc_hd__a21o_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$400 U$$948/A1 U$$278/X U$$539/A1 U$$279/X VGND VGND VPWR VPWR U$$401/A sky130_fd_sc_hd__a22o_1
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_633_ _633_/CLK _633_/D VGND VGND VPWR VPWR _633_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$411 _621_/Q VGND VGND VPWR VPWR U$$411/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$583 final_adder.U$$710/A final_adder.U$$710/B final_adder.U$$583/B1
+ VGND VGND VPWR VPWR final_adder.U$$711/B sky130_fd_sc_hd__a21o_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$422 U$$422/A U$$530/B VGND VGND VPWR VPWR U$$422/X sky130_fd_sc_hd__xor2_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_35_3 dadda_fa_3_35_3/A dadda_fa_3_35_3/B dadda_fa_3_35_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/B dadda_fa_4_35_2/CIN sky130_fd_sc_hd__fa_1
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$433 _559_/Q U$$491/A2 U$$983/A1 U$$416/X VGND VGND VPWR VPWR U$$434/A sky130_fd_sc_hd__a22o_1
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$444 U$$444/A U$$530/B VGND VGND VPWR VPWR U$$444/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_83_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _633_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$455 _570_/Q U$$491/A2 U$$46/A1 U$$416/X VGND VGND VPWR VPWR U$$456/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_28_2 dadda_fa_3_28_2/A dadda_fa_3_28_2/B dadda_fa_3_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/A dadda_fa_4_28_2/B sky130_fd_sc_hd__fa_1
XFILLER_45_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_564_ _637_/CLK _564_/D VGND VGND VPWR VPWR _564_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$466 U$$466/A _623_/Q VGND VGND VPWR VPWR U$$466/X sky130_fd_sc_hd__xor2_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$477 U$$66/A1 U$$491/A2 U$$68/A1 U$$416/X VGND VGND VPWR VPWR U$$478/A sky130_fd_sc_hd__a22o_1
XU$$488 U$$488/A U$$530/B VGND VGND VPWR VPWR U$$488/X sky130_fd_sc_hd__xor2_1
XFILLER_72_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$499 U$$771/B1 U$$545/A2 U$$90/A1 U$$416/X VGND VGND VPWR VPWR U$$500/A sky130_fd_sc_hd__a22o_1
XFILLER_60_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_495_ _495_/CLK _495_/D VGND VGND VPWR VPWR _495_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_2_31_4 U$$1665/X U$$1798/X VGND VGND VPWR VPWR dadda_fa_3_32_2/A dadda_fa_4_31_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_7_1_0 U$$9/X input168/X VGND VGND VPWR VPWR _426_/D _297_/D sky130_fd_sc_hd__ha_1
XFILLER_78_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk _560_/CLK VGND VGND VPWR VPWR _645_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_30_2 U$$865/X U$$998/X U$$1131/X VGND VGND VPWR VPWR dadda_fa_3_31_1/CIN
+ dadda_fa_3_30_3/B sky130_fd_sc_hd__fa_1
XFILLER_39_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1150 U$$54/A1 U$$1200/A2 U$$56/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1151/A sky130_fd_sc_hd__a22o_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1161 U$$1161/A U$$1167/B VGND VGND VPWR VPWR U$$1161/X sky130_fd_sc_hd__xor2_1
XU$$1172 U$$2953/A1 U$$1218/A2 U$$76/B1 U$$1218/B2 VGND VGND VPWR VPWR U$$1173/A sky130_fd_sc_hd__a22o_1
XFILLER_149_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1183 U$$1183/A U$$1232/A VGND VGND VPWR VPWR U$$1183/X sky130_fd_sc_hd__xor2_1
XU$$1194 U$$96/B1 U$$1218/A2 U$$785/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1195/A sky130_fd_sc_hd__a22o_1
XFILLER_31_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_753__805 VGND VGND VPWR VPWR _753__805/HI U$$3696/B1 sky130_fd_sc_hd__conb_1
XFILLER_176_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_82_5 U$$3230/X U$$3363/X U$$3496/X VGND VGND VPWR VPWR dadda_fa_2_83_3/A
+ dadda_fa_2_82_5/B sky130_fd_sc_hd__fa_1
XFILLER_160_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_75_4 U$$3216/X U$$3349/X U$$3482/X VGND VGND VPWR VPWR dadda_fa_2_76_1/CIN
+ dadda_fa_2_75_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_3 U$$3734/X U$$3867/X U$$4000/X VGND VGND VPWR VPWR dadda_fa_2_69_1/B
+ dadda_fa_2_68_4/B sky130_fd_sc_hd__fa_2
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_45_2 dadda_fa_4_45_2/A dadda_fa_4_45_2/B dadda_fa_4_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/CIN dadda_fa_5_45_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_38_1 dadda_fa_4_38_1/A dadda_fa_4_38_1/B dadda_fa_4_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/B dadda_fa_5_38_1/B sky130_fd_sc_hd__fa_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_65_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _573_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_7_15_0 dadda_fa_7_15_0/A dadda_fa_7_15_0/B dadda_fa_7_15_0/CIN VGND VGND
+ VPWR VPWR _440_/D _311_/D sky130_fd_sc_hd__fa_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ _280_/CLK _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_70_3 U$$1610/X U$$1743/X U$$1876/X VGND VGND VPWR VPWR dadda_fa_1_71_7/B
+ dadda_fa_1_70_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_63_2 U$$931/X U$$1064/X U$$1197/X VGND VGND VPWR VPWR dadda_fa_1_64_6/A
+ dadda_fa_1_63_8/A sky130_fd_sc_hd__fa_1
XFILLER_65_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_1 dadda_fa_3_40_1/A dadda_fa_3_40_1/B dadda_fa_3_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/CIN dadda_fa_4_40_2/A sky130_fd_sc_hd__fa_2
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_1 U$$518/X U$$651/X U$$784/X VGND VGND VPWR VPWR dadda_fa_1_57_7/CIN
+ dadda_fa_1_56_8/CIN sky130_fd_sc_hd__fa_2
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk _536_/CLK VGND VGND VPWR VPWR _597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_33_0 input183/X dadda_fa_3_33_0/B dadda_fa_3_33_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_34_0/B dadda_fa_4_33_1/CIN sky130_fd_sc_hd__fa_2
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$230 U$$230/A U$$242/B VGND VGND VPWR VPWR U$$230/X sky130_fd_sc_hd__xor2_1
XFILLER_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$391 final_adder.U$$354/B final_adder.U$$638/B final_adder.U$$325/X
+ VGND VGND VPWR VPWR final_adder.U$$646/B sky130_fd_sc_hd__a21o_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _622_/CLK _616_/D VGND VGND VPWR VPWR U$$1/A sky130_fd_sc_hd__dfxtp_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$241 U$$926/A1 U$$141/X U$$928/A1 U$$142/X VGND VGND VPWR VPWR U$$242/A sky130_fd_sc_hd__a22o_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$252 U$$252/A U$$274/A VGND VGND VPWR VPWR U$$252/X sky130_fd_sc_hd__xor2_1
XFILLER_18_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$263 U$$948/A1 U$$141/X U$$950/A1 U$$142/X VGND VGND VPWR VPWR U$$264/A sky130_fd_sc_hd__a22o_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$274 U$$274/A VGND VGND VPWR VPWR U$$274/Y sky130_fd_sc_hd__inv_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$285 U$$285/A U$$357/B VGND VGND VPWR VPWR U$$285/X sky130_fd_sc_hd__xor2_1
X_547_ _678_/CLK _547_/D VGND VGND VPWR VPWR _547_/Q sky130_fd_sc_hd__dfxtp_2
XU$$296 U$$979/B1 U$$278/X U$$983/A1 U$$279/X VGND VGND VPWR VPWR U$$297/A sky130_fd_sc_hd__a22o_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_478_ _480_/CLK _478_/D VGND VGND VPWR VPWR _478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2 U$$3/A VGND VGND VPWR VPWR U$$2/Y sky130_fd_sc_hd__inv_1
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput305 _196_/Q VGND VGND VPWR VPWR o[28] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_4 input248/X dadda_fa_2_92_4/B dadda_fa_2_92_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_93_1/CIN dadda_fa_3_92_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput316 _206_/Q VGND VGND VPWR VPWR o[38] sky130_fd_sc_hd__buf_2
Xoutput327 _216_/Q VGND VGND VPWR VPWR o[48] sky130_fd_sc_hd__buf_2
XFILLER_142_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput338 _226_/Q VGND VGND VPWR VPWR o[58] sky130_fd_sc_hd__buf_2
XFILLER_99_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput349 _236_/Q VGND VGND VPWR VPWR o[68] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_3 dadda_fa_2_85_3/A dadda_fa_2_85_3/B dadda_fa_2_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/B dadda_fa_3_85_3/B sky130_fd_sc_hd__fa_2
XFILLER_114_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_78_2 dadda_fa_2_78_2/A dadda_fa_2_78_2/B dadda_fa_2_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/A dadda_fa_3_78_3/A sky130_fd_sc_hd__fa_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_55_1 dadda_fa_5_55_1/A dadda_fa_5_55_1/B dadda_fa_5_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/B dadda_fa_7_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_171_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_48_0 dadda_fa_5_48_0/A dadda_fa_5_48_0/B dadda_fa_5_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/A dadda_fa_6_48_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_2_22_0 U$$51/X U$$184/X VGND VGND VPWR VPWR dadda_fa_3_23_3/CIN dadda_fa_4_22_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_clk _536_/CLK VGND VGND VPWR VPWR _612_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_101_1 U$$3002/X U$$3135/X U$$3268/X VGND VGND VPWR VPWR dadda_fa_3_102_2/A
+ dadda_fa_3_101_3/B sky130_fd_sc_hd__fa_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_122_0 U$$4241/X U$$4374/X U$$4507/X VGND VGND VPWR VPWR dadda_fa_6_123_0/A
+ dadda_fa_6_122_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_80_2 U$$1896/X U$$2029/X U$$2162/X VGND VGND VPWR VPWR dadda_fa_2_81_1/B
+ dadda_fa_2_80_4/A sky130_fd_sc_hd__fa_1
XFILLER_104_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_73_1 U$$2281/X U$$2414/X U$$2547/X VGND VGND VPWR VPWR dadda_fa_2_74_0/CIN
+ dadda_fa_2_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_50_0 dadda_fa_4_50_0/A dadda_fa_4_50_0/B dadda_fa_4_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/A dadda_fa_5_50_1/A sky130_fd_sc_hd__fa_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_66_0 U$$2533/X U$$2666/X U$$2799/X VGND VGND VPWR VPWR dadda_fa_2_67_0/B
+ dadda_fa_2_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_150_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_38_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _500_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2609 U$$2609/A1 U$$2729/A2 U$$8/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2610/A sky130_fd_sc_hd__a22o_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1908 U$$1908/A _643_/Q VGND VGND VPWR VPWR U$$1908/X sky130_fd_sc_hd__xor2_1
X_401_ _535_/CLK _401_/D VGND VGND VPWR VPWR _401_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1919 _644_/Q VGND VGND VPWR VPWR U$$1921/B sky130_fd_sc_hd__inv_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_332_ _333_/CLK _332_/D VGND VGND VPWR VPWR _332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_263_ _267_/CLK _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_1
X_194_ _329_/CLK _194_/D VGND VGND VPWR VPWR _194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_95_2 dadda_fa_3_95_2/A dadda_fa_3_95_2/B dadda_fa_3_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/A dadda_fa_4_95_2/B sky130_fd_sc_hd__fa_2
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_88_1 dadda_fa_3_88_1/A dadda_fa_3_88_1/B dadda_fa_3_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/CIN dadda_fa_4_88_2/A sky130_fd_sc_hd__fa_2
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_65_0 dadda_fa_6_65_0/A dadda_fa_6_65_0/B dadda_fa_6_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_66_0/B dadda_fa_7_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4501 U$$4501/A U$$4501/B VGND VGND VPWR VPWR U$$4501/X sky130_fd_sc_hd__xor2_1
XU$$4512 U$$539/A1 U$$4388/X U$$4514/A1 U$$4389/X VGND VGND VPWR VPWR U$$4513/A sky130_fd_sc_hd__a22o_1
XU$$3800 U$$3800/A _671_/Q VGND VGND VPWR VPWR U$$3800/X sky130_fd_sc_hd__xor2_1
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$15 U$$15/A U$$9/B VGND VGND VPWR VPWR U$$15/X sky130_fd_sc_hd__xor2_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$26 U$$26/A1 U$$4/X U$$28/A1 U$$5/X VGND VGND VPWR VPWR U$$27/A sky130_fd_sc_hd__a22o_1
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3811 U$$934/A1 U$$3703/X _605_/Q U$$3704/X VGND VGND VPWR VPWR U$$3812/A sky130_fd_sc_hd__a22o_1
XU$$37 U$$37/A U$$3/A VGND VGND VPWR VPWR U$$37/X sky130_fd_sc_hd__xor2_1
XU$$3822 U$$3822/A U$$3835/A VGND VGND VPWR VPWR U$$3822/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_1 U$$4098/X U$$4231/X U$$4364/X VGND VGND VPWR VPWR dadda_fa_5_118_0/B
+ dadda_fa_5_117_1/B sky130_fd_sc_hd__fa_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk _369_/CLK VGND VGND VPWR VPWR _492_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3833 U$$819/A1 U$$3703/X U$$3833/B1 U$$3704/X VGND VGND VPWR VPWR U$$3834/A sky130_fd_sc_hd__a22o_1
XFILLER_64_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3844 U$$4255/A1 U$$3912/A2 U$$969/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3845/A
+ sky130_fd_sc_hd__a22o_1
XU$$48 U$$48/A1 U$$4/X U$$50/A1 U$$5/X VGND VGND VPWR VPWR U$$49/A sky130_fd_sc_hd__a22o_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$59 U$$59/A U$$3/A VGND VGND VPWR VPWR U$$59/X sky130_fd_sc_hd__xor2_1
XU$$3855 U$$3855/A U$$3929/B VGND VGND VPWR VPWR U$$3855/X sky130_fd_sc_hd__xor2_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3866 _563_/Q U$$3912/A2 _564_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3867/A sky130_fd_sc_hd__a22o_1
XFILLER_18_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3877 U$$3877/A U$$3893/B VGND VGND VPWR VPWR U$$3877/X sky130_fd_sc_hd__xor2_1
XFILLER_75_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3888 U$$52/A1 U$$3912/A2 U$$4438/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3889/A sky130_fd_sc_hd__a22o_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3899 U$$3899/A U$$3969/B VGND VGND VPWR VPWR U$$3899/X sky130_fd_sc_hd__xor2_1
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_90_1 U$$3645/X U$$3778/X U$$3911/X VGND VGND VPWR VPWR dadda_fa_3_91_0/CIN
+ dadda_fa_3_90_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_173_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_83_0 U$$4163/X U$$4296/X U$$4429/X VGND VGND VPWR VPWR dadda_fa_3_84_0/B
+ dadda_fa_3_83_2/B sky130_fd_sc_hd__fa_2
XFILLER_82_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_52_6 U$$2771/X U$$2904/X U$$3037/X VGND VGND VPWR VPWR dadda_fa_2_53_2/B
+ dadda_fa_2_52_5/B sky130_fd_sc_hd__fa_2
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_4_0 dadda_fa_7_4_0/A dadda_fa_7_4_0/B dadda_fa_7_4_0/CIN VGND VGND VPWR
+ VPWR _429_/D _300_/D sky130_fd_sc_hd__fa_1
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_759__811 VGND VGND VPWR VPWR _759__811/HI U$$4/A3 sky130_fd_sc_hd__conb_1
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_82_0 dadda_fa_7_82_0/A dadda_fa_7_82_0/B dadda_fa_7_82_0/CIN VGND VGND
+ VPWR VPWR _507_/D _378_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_98_0 dadda_fa_4_98_0/A dadda_fa_4_98_0/B dadda_fa_4_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/A dadda_fa_5_98_1/A sky130_fd_sc_hd__fa_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3107 U$$3107/A _661_/Q VGND VGND VPWR VPWR U$$3107/X sky130_fd_sc_hd__xor2_1
XFILLER_47_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3118 U$$787/B1 U$$3018/X U$$654/A1 U$$3019/X VGND VGND VPWR VPWR U$$3119/A sky130_fd_sc_hd__a22o_1
XU$$3129 U$$3129/A U$$3129/B VGND VGND VPWR VPWR U$$3129/X sky130_fd_sc_hd__xor2_1
XFILLER_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2406 U$$2406/A U$$2432/B VGND VGND VPWR VPWR U$$2406/X sky130_fd_sc_hd__xor2_1
XU$$2417 U$$4335/A1 U$$2421/A2 _593_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2418/A sky130_fd_sc_hd__a22o_1
XFILLER_74_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2428 U$$2428/A U$$2464/B VGND VGND VPWR VPWR U$$2428/X sky130_fd_sc_hd__xor2_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2439 U$$4494/A1 U$$2463/A2 U$$4496/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2440/A
+ sky130_fd_sc_hd__a22o_1
XU$$1705 U$$1705/A U$$1739/B VGND VGND VPWR VPWR U$$1705/X sky130_fd_sc_hd__xor2_1
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1716 U$$892/B1 U$$1726/A2 U$$74/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1717/A sky130_fd_sc_hd__a22o_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1727 U$$1727/A U$$1727/B VGND VGND VPWR VPWR U$$1727/X sky130_fd_sc_hd__xor2_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1738 U$$92/B1 U$$1770/A2 U$$96/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1739/A sky130_fd_sc_hd__a22o_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1749 U$$1749/A _641_/Q VGND VGND VPWR VPWR U$$1749/X sky130_fd_sc_hd__xor2_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _452_/CLK _315_/D VGND VGND VPWR VPWR _315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_246_ _501_/CLK _246_/D VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 a[22] VGND VGND VPWR VPWR _638_/D sky130_fd_sc_hd__buf_2
XFILLER_11_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput26 a[32] VGND VGND VPWR VPWR _648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput37 a[42] VGND VGND VPWR VPWR _658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput48 a[52] VGND VGND VPWR VPWR _668_/D sky130_fd_sc_hd__clkbuf_1
Xinput59 a[62] VGND VGND VPWR VPWR _678_/D sky130_fd_sc_hd__clkbuf_1
X_177_ _462_/CLK _177_/D VGND VGND VPWR VPWR _177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_62_5 dadda_fa_2_62_5/A dadda_fa_2_62_5/B dadda_fa_2_62_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_2/A dadda_fa_4_62_0/A sky130_fd_sc_hd__fa_2
Xrepeater605 _621_/Q VGND VGND VPWR VPWR U$$391/B sky130_fd_sc_hd__buf_12
XFILLER_111_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater616 U$$4514/A1 VGND VGND VPWR VPWR U$$952/A1 sky130_fd_sc_hd__buf_12
XFILLER_96_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater627 _608_/Q VGND VGND VPWR VPWR U$$4504/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_55_4 dadda_fa_2_55_4/A dadda_fa_2_55_4/B dadda_fa_2_55_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/CIN dadda_fa_3_55_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_38_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater638 U$$4492/A1 VGND VGND VPWR VPWR U$$930/A1 sky130_fd_sc_hd__buf_12
Xrepeater649 _598_/Q VGND VGND VPWR VPWR U$$4484/A1 sky130_fd_sc_hd__buf_12
XU$$4320 U$$4320/A U$$4332/B VGND VGND VPWR VPWR U$$4320/X sky130_fd_sc_hd__xor2_1
XU$$4331 U$$632/A1 U$$4251/X U$$771/A1 U$$4252/X VGND VGND VPWR VPWR U$$4332/A sky130_fd_sc_hd__a22o_1
XFILLER_93_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4342 U$$4342/A U$$4384/A VGND VGND VPWR VPWR U$$4342/X sky130_fd_sc_hd__xor2_2
XU$$4353 U$$654/A1 U$$4377/A2 U$$4492/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4354/A
+ sky130_fd_sc_hd__a22o_1
XU$$4364 U$$4364/A U$$4384/A VGND VGND VPWR VPWR U$$4364/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_3 dadda_fa_2_48_3/A dadda_fa_2_48_3/B dadda_fa_2_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/B dadda_fa_3_48_3/B sky130_fd_sc_hd__fa_1
XU$$3630 U$$4178/A1 U$$3668/A2 _583_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3631/A sky130_fd_sc_hd__a22o_1
XU$$4375 U$$539/A1 U$$4377/A2 _613_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4376/A sky130_fd_sc_hd__a22o_1
XU$$3641 U$$3641/A U$$3699/A VGND VGND VPWR VPWR U$$3641/X sky130_fd_sc_hd__xor2_1
XU$$4386 U$$4386/A VGND VGND VPWR VPWR U$$4386/Y sky130_fd_sc_hd__inv_1
XFILLER_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4397 U$$4397/A U$$4397/B VGND VGND VPWR VPWR U$$4397/X sky130_fd_sc_hd__xor2_2
XU$$3652 U$$90/A1 U$$3566/X U$$4476/A1 U$$3567/X VGND VGND VPWR VPWR U$$3653/A sky130_fd_sc_hd__a22o_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3663 U$$3663/A U$$3699/A VGND VGND VPWR VPWR U$$3663/X sky130_fd_sc_hd__xor2_1
XU$$3674 U$$4496/A1 U$$3566/X _605_/Q U$$3567/X VGND VGND VPWR VPWR U$$3675/A sky130_fd_sc_hd__a22o_1
XU$$2940 U$$2940/A U$$2960/B VGND VGND VPWR VPWR U$$2940/X sky130_fd_sc_hd__xor2_1
XU$$3685 U$$3685/A U$$3698/A VGND VGND VPWR VPWR U$$3685/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_18_1 dadda_fa_5_18_1/A dadda_fa_5_18_1/B dadda_fa_5_18_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/B dadda_fa_7_18_0/A sky130_fd_sc_hd__fa_1
XFILLER_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3696 U$$819/A1 U$$3566/X U$$3696/B1 U$$3567/X VGND VGND VPWR VPWR U$$3697/A sky130_fd_sc_hd__a22o_1
XFILLER_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2951 U$$4045/B1 U$$2975/A2 U$$2953/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2952/A
+ sky130_fd_sc_hd__a22o_1
XU$$2962 U$$2962/A _659_/Q VGND VGND VPWR VPWR U$$2962/X sky130_fd_sc_hd__xor2_1
XU$$2973 U$$94/B1 U$$3009/A2 U$$98/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2974/A sky130_fd_sc_hd__a22o_1
XU$$2984 U$$2984/A U$$3004/B VGND VGND VPWR VPWR U$$2984/X sky130_fd_sc_hd__xor2_1
XU$$2995 U$$940/A1 U$$3009/A2 U$$942/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2996/A sky130_fd_sc_hd__a22o_1
XFILLER_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_clk _431_/CLK VGND VGND VPWR VPWR _425_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_50_3 U$$1304/X U$$1437/X U$$1570/X VGND VGND VPWR VPWR dadda_fa_2_51_1/B
+ dadda_fa_2_50_4/B sky130_fd_sc_hd__fa_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$807 U$$944/A1 U$$817/A2 U$$946/A1 U$$817/B2 VGND VGND VPWR VPWR U$$808/A sky130_fd_sc_hd__a22o_1
XFILLER_84_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$818 U$$818/A _627_/Q VGND VGND VPWR VPWR U$$818/X sky130_fd_sc_hd__xor2_1
XFILLER_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_43_2 U$$891/X U$$1024/X U$$1157/X VGND VGND VPWR VPWR dadda_fa_2_44_3/B
+ dadda_fa_2_43_5/B sky130_fd_sc_hd__fa_1
XU$$829 U$$829/A U$$903/B VGND VGND VPWR VPWR U$$829/X sky130_fd_sc_hd__xor2_2
Xdadda_fa_4_20_1 dadda_fa_4_20_1/A dadda_fa_4_20_1/B dadda_fa_4_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/B dadda_fa_5_20_1/B sky130_fd_sc_hd__fa_2
XFILLER_25_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_13_0 U$$33/X U$$166/X U$$299/X VGND VGND VPWR VPWR dadda_fa_5_14_0/A dadda_fa_5_13_1/A
+ sky130_fd_sc_hd__fa_2
XFILLER_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_65_3 dadda_fa_3_65_3/A dadda_fa_3_65_3/B dadda_fa_3_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/B dadda_fa_4_65_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_58_2 dadda_fa_3_58_2/A dadda_fa_3_58_2/B dadda_fa_3_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/A dadda_fa_4_58_2/B sky130_fd_sc_hd__fa_1
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_28_0 dadda_fa_6_28_0/A dadda_fa_6_28_0/B dadda_fa_6_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_29_0/B dadda_fa_7_28_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2203 U$$2203/A U$$2257/B VGND VGND VPWR VPWR U$$2203/X sky130_fd_sc_hd__xor2_1
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2214 U$$979/B1 U$$2270/A2 U$$983/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2215/A sky130_fd_sc_hd__a22o_1
XU$$2225 U$$2225/A U$$2257/B VGND VGND VPWR VPWR U$$2225/X sky130_fd_sc_hd__xor2_1
XU$$2236 U$$4289/B1 U$$2270/A2 U$$4291/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2237/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1502 U$$952/B1 U$$1374/X U$$956/A1 U$$1375/X VGND VGND VPWR VPWR U$$1503/A sky130_fd_sc_hd__a22o_1
XU$$2247 U$$2247/A U$$2257/B VGND VGND VPWR VPWR U$$2247/X sky130_fd_sc_hd__xor2_1
XFILLER_16_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1513 U$$1513/A1 U$$1511/X U$$8/A1 U$$1512/X VGND VGND VPWR VPWR U$$1514/A sky130_fd_sc_hd__a22o_1
XU$$2258 U$$3489/B1 U$$2316/A2 U$$68/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2259/A sky130_fd_sc_hd__a22o_1
XU$$2269 U$$2269/A U$$2327/B VGND VGND VPWR VPWR U$$2269/X sky130_fd_sc_hd__xor2_1
XU$$1524 U$$1524/A U$$1580/B VGND VGND VPWR VPWR U$$1524/X sky130_fd_sc_hd__xor2_1
XU$$1535 U$$987/A1 U$$1591/A2 U$$28/B1 U$$1591/B2 VGND VGND VPWR VPWR U$$1536/A sky130_fd_sc_hd__a22o_1
XFILLER_43_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1546 U$$1546/A U$$1580/B VGND VGND VPWR VPWR U$$1546/X sky130_fd_sc_hd__xor2_1
XU$$1557 U$$50/A1 U$$1605/A2 U$$2790/B1 U$$1605/B2 VGND VGND VPWR VPWR U$$1558/A sky130_fd_sc_hd__a22o_1
XFILLER_31_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1568 U$$1568/A U$$1614/B VGND VGND VPWR VPWR U$$1568/X sky130_fd_sc_hd__xor2_1
XU$$1579 U$$892/B1 U$$1605/A2 U$$74/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1580/A sky130_fd_sc_hd__a22o_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_229_ _499_/CLK _229_/D VGND VGND VPWR VPWR _229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_2 dadda_fa_2_60_2/A dadda_fa_2_60_2/B dadda_fa_2_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/A dadda_fa_3_60_3/A sky130_fd_sc_hd__fa_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater402 U$$3840/X VGND VGND VPWR VPWR U$$3970/A2 sky130_fd_sc_hd__buf_12
XFILLER_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$209 final_adder.U$$703/A final_adder.U$$575/B1 final_adder.U$$209/B1
+ VGND VGND VPWR VPWR final_adder.U$$209/X sky130_fd_sc_hd__a21o_1
Xrepeater413 U$$3155/X VGND VGND VPWR VPWR U$$3241/A2 sky130_fd_sc_hd__buf_12
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater424 U$$2574/A2 VGND VGND VPWR VPWR U$$2584/A2 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_53_1 dadda_fa_2_53_1/A dadda_fa_2_53_1/B dadda_fa_2_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/CIN dadda_fa_3_53_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater435 U$$2052/A2 VGND VGND VPWR VPWR U$$2048/A2 sky130_fd_sc_hd__buf_12
XFILLER_66_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater446 U$$1474/A2 VGND VGND VPWR VPWR U$$1472/A2 sky130_fd_sc_hd__buf_12
Xrepeater457 U$$817/B2 VGND VGND VPWR VPWR U$$785/B2 sky130_fd_sc_hd__buf_12
Xdadda_fa_5_30_0 dadda_fa_5_30_0/A dadda_fa_5_30_0/B dadda_fa_5_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/A dadda_fa_6_30_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater468 U$$3704/X VGND VGND VPWR VPWR U$$3795/B2 sky130_fd_sc_hd__buf_12
XU$$4150 U$$4424/A1 U$$4114/X U$$4289/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4151/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_0 U$$2759/X U$$2892/X U$$3025/X VGND VGND VPWR VPWR dadda_fa_3_47_0/B
+ dadda_fa_3_46_2/B sky130_fd_sc_hd__fa_1
Xrepeater479 U$$3019/X VGND VGND VPWR VPWR U$$3146/B2 sky130_fd_sc_hd__buf_12
XU$$4161 U$$4161/A U$$4247/A VGND VGND VPWR VPWR U$$4161/X sky130_fd_sc_hd__xor2_1
XFILLER_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4172 U$$4446/A1 U$$4114/X _580_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4173/A sky130_fd_sc_hd__a22o_1
XFILLER_26_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4183 U$$4183/A U$$4246/A VGND VGND VPWR VPWR U$$4183/X sky130_fd_sc_hd__xor2_1
XFILLER_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4194 U$$632/A1 U$$4198/A2 U$$771/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4195/A sky130_fd_sc_hd__a22o_1
XU$$3460 U$$3460/A U$$3561/A VGND VGND VPWR VPWR U$$3460/X sky130_fd_sc_hd__xor2_1
XFILLER_81_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3471 U$$4291/B1 U$$3525/A2 U$$4156/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3472/A
+ sky130_fd_sc_hd__a22o_1
XU$$3482 U$$3482/A U$$3496/B VGND VGND VPWR VPWR U$$3482/X sky130_fd_sc_hd__xor2_1
XU$$3493 U$$4178/A1 U$$3525/A2 U$$892/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3494/A
+ sky130_fd_sc_hd__a22o_1
XU$$2770 _563_/Q U$$2796/A2 _564_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2771/A sky130_fd_sc_hd__a22o_1
XU$$2781 U$$2781/A U$$2839/B VGND VGND VPWR VPWR U$$2781/X sky130_fd_sc_hd__xor2_1
X_721__773 VGND VGND VPWR VPWR _721__773/HI U$$1641/B1 sky130_fd_sc_hd__conb_1
XU$$2792 U$$50/B1 U$$2796/A2 U$$876/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2793/A sky130_fd_sc_hd__a22o_1
XFILLER_178_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_75_2 dadda_fa_4_75_2/A dadda_fa_4_75_2/B dadda_fa_4_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/CIN dadda_fa_5_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_68_1 dadda_fa_4_68_1/A dadda_fa_4_68_1/B dadda_fa_4_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/B dadda_fa_5_68_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput205 c[53] VGND VGND VPWR VPWR input205/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput216 c[63] VGND VGND VPWR VPWR input216/X sky130_fd_sc_hd__buf_2
Xdadda_fa_7_45_0 dadda_fa_7_45_0/A dadda_fa_7_45_0/B dadda_fa_7_45_0/CIN VGND VGND
+ VPWR VPWR _470_/D _341_/D sky130_fd_sc_hd__fa_2
Xinput227 c[73] VGND VGND VPWR VPWR input227/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput238 c[83] VGND VGND VPWR VPWR input238/X sky130_fd_sc_hd__buf_2
Xdadda_ha_1_35_0 U$$77/X U$$210/X VGND VGND VPWR VPWR dadda_fa_2_36_5/B dadda_fa_3_35_0/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$710 final_adder.U$$710/A final_adder.U$$710/B VGND VGND VPWR VPWR
+ _256_/D sky130_fd_sc_hd__xor2_1
Xinput249 c[93] VGND VGND VPWR VPWR input249/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$721 final_adder.U$$721/A final_adder.U$$721/B VGND VGND VPWR VPWR
+ _267_/D sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$732 final_adder.U$$732/A final_adder.U$$732/B VGND VGND VPWR VPWR
+ _278_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$743 final_adder.U$$743/A final_adder.U$$743/B VGND VGND VPWR VPWR
+ _289_/D sky130_fd_sc_hd__xor2_1
XU$$604 U$$878/A1 U$$682/A2 U$$58/A1 U$$553/X VGND VGND VPWR VPWR U$$605/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$615 U$$615/A _625_/Q VGND VGND VPWR VPWR U$$615/X sky130_fd_sc_hd__xor2_1
X_580_ _581_/CLK _580_/D VGND VGND VPWR VPWR _580_/Q sky130_fd_sc_hd__dfxtp_4
XU$$626 U$$78/A1 U$$626/A2 U$$80/A1 U$$553/X VGND VGND VPWR VPWR U$$627/A sky130_fd_sc_hd__a22o_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$637 U$$637/A U$$661/B VGND VGND VPWR VPWR U$$637/X sky130_fd_sc_hd__xor2_1
XFILLER_84_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$648 U$$785/A1 U$$682/A2 U$$924/A1 U$$553/X VGND VGND VPWR VPWR U$$649/A sky130_fd_sc_hd__a22o_1
XU$$659 U$$659/A U$$661/B VGND VGND VPWR VPWR U$$659/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_70_1 dadda_fa_3_70_1/A dadda_fa_3_70_1/B dadda_fa_3_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/CIN dadda_fa_4_70_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_63_0 dadda_fa_3_63_0/A dadda_fa_3_63_0/B dadda_fa_3_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/B dadda_fa_4_63_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2000 U$$82/A1 U$$2052/A2 U$$632/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2001/A sky130_fd_sc_hd__a22o_1
XU$$2011 U$$2011/A U$$2023/B VGND VGND VPWR VPWR U$$2011/X sky130_fd_sc_hd__xor2_1
XU$$2022 U$$926/A1 U$$2036/A2 U$$928/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$2023/A sky130_fd_sc_hd__a22o_1
XFILLER_35_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2033 U$$2033/A U$$2055/A VGND VGND VPWR VPWR U$$2033/X sky130_fd_sc_hd__xor2_1
XU$$2044 U$$948/A1 U$$2052/A2 U$$950/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2045/A sky130_fd_sc_hd__a22o_1
XU$$1310 U$$1310/A U$$1369/A VGND VGND VPWR VPWR U$$1310/X sky130_fd_sc_hd__xor2_1
XU$$2055 U$$2055/A VGND VGND VPWR VPWR U$$2055/Y sky130_fd_sc_hd__inv_1
XFILLER_90_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2066 U$$2066/A U$$2186/B VGND VGND VPWR VPWR U$$2066/X sky130_fd_sc_hd__xor2_1
XU$$1321 U$$88/A1 U$$1367/A2 U$$912/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1322/A sky130_fd_sc_hd__a22o_1
XU$$1332 U$$1332/A U$$1336/B VGND VGND VPWR VPWR U$$1332/X sky130_fd_sc_hd__xor2_1
XU$$2077 U$$22/A1 U$$2059/X _560_/Q U$$2117/B2 VGND VGND VPWR VPWR U$$2078/A sky130_fd_sc_hd__a22o_1
XU$$2088 U$$2088/A U$$2118/B VGND VGND VPWR VPWR U$$2088/X sky130_fd_sc_hd__xor2_1
XU$$1343 _603_/Q U$$1367/A2 U$$934/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1344/A sky130_fd_sc_hd__a22o_1
XU$$1354 U$$1354/A U$$1369/A VGND VGND VPWR VPWR U$$1354/X sky130_fd_sc_hd__xor2_1
XU$$2099 U$$4291/A1 U$$2117/A2 U$$868/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2100/A
+ sky130_fd_sc_hd__a22o_1
XU$$1365 _614_/Q U$$1367/A2 _615_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1366/A sky130_fd_sc_hd__a22o_1
XU$$1376 U$$1376/A1 U$$1474/A2 U$$8/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1377/A sky130_fd_sc_hd__a22o_1
XU$$1387 U$$1387/A U$$1479/B VGND VGND VPWR VPWR U$$1387/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_120_0 dadda_fa_7_120_0/A dadda_fa_7_120_0/B dadda_fa_7_120_0/CIN VGND
+ VGND VPWR VPWR _545_/D _416_/D sky130_fd_sc_hd__fa_2
XU$$1398 U$$987/A1 U$$1474/A2 U$$28/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1399/A sky130_fd_sc_hd__a22o_1
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_85_1 dadda_fa_5_85_1/A dadda_fa_5_85_1/B dadda_fa_5_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/B dadda_fa_7_85_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_78_0 dadda_fa_5_78_0/A dadda_fa_5_78_0/B dadda_fa_5_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/A dadda_fa_6_78_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_77_8 input231/X dadda_fa_1_77_8/B dadda_fa_1_77_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_78_3/A dadda_fa_3_77_0/A sky130_fd_sc_hd__fa_2
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$50 _474_/Q _346_/Q VGND VGND VPWR VPWR final_adder.U$$545/B1 final_adder.U$$672/A
+ sky130_fd_sc_hd__ha_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$61 _485_/Q _357_/Q VGND VGND VPWR VPWR final_adder.U$$189/B1 final_adder.U$$683/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3290 _665_/Q VGND VGND VPWR VPWR U$$3290/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$72 _496_/Q _368_/Q VGND VGND VPWR VPWR final_adder.U$$567/B1 final_adder.U$$694/A
+ sky130_fd_sc_hd__ha_2
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$83 _507_/Q _379_/Q VGND VGND VPWR VPWR final_adder.U$$211/B1 final_adder.U$$705/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$94 _518_/Q _390_/Q VGND VGND VPWR VPWR final_adder.U$$589/B1 final_adder.U$$716/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_80_0 dadda_fa_4_80_0/A dadda_fa_4_80_0/B dadda_fa_4_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/A dadda_fa_5_80_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_101_3 dadda_fa_3_101_3/A dadda_fa_3_101_3/B dadda_fa_3_101_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/B dadda_fa_4_101_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$551 final_adder.U$$678/A final_adder.U$$678/B final_adder.U$$551/B1
+ VGND VGND VPWR VPWR final_adder.U$$679/B sky130_fd_sc_hd__a21o_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_632_ _632_/CLK _632_/D VGND VGND VPWR VPWR _632_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$401 U$$401/A _621_/Q VGND VGND VPWR VPWR U$$401/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_108_0 dadda_fa_6_108_0/A dadda_fa_6_108_0/B dadda_fa_6_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_109_0/B dadda_fa_7_108_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$573 final_adder.U$$700/A final_adder.U$$700/B final_adder.U$$573/B1
+ VGND VGND VPWR VPWR final_adder.U$$701/B sky130_fd_sc_hd__a21o_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$412 _622_/Q VGND VGND VPWR VPWR U$$414/B sky130_fd_sc_hd__inv_1
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$423 U$$971/A1 U$$491/A2 U$$12/B1 U$$416/X VGND VGND VPWR VPWR U$$424/A sky130_fd_sc_hd__a22o_1
XFILLER_91_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$595 final_adder.U$$722/A final_adder.U$$722/B final_adder.U$$595/B1
+ VGND VGND VPWR VPWR final_adder.U$$723/B sky130_fd_sc_hd__a21o_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$434 U$$434/A U$$530/B VGND VGND VPWR VPWR U$$434/X sky130_fd_sc_hd__xor2_1
XFILLER_72_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$445 U$$34/A1 U$$545/A2 U$$36/A1 U$$416/X VGND VGND VPWR VPWR U$$446/A sky130_fd_sc_hd__a22o_1
X_563_ _637_/CLK _563_/D VGND VGND VPWR VPWR _563_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$456 U$$456/A U$$530/B VGND VGND VPWR VPWR U$$456/X sky130_fd_sc_hd__xor2_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_3 dadda_fa_3_28_3/A dadda_fa_3_28_3/B dadda_fa_3_28_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/B dadda_fa_4_28_2/CIN sky130_fd_sc_hd__fa_2
XU$$467 U$$878/A1 U$$491/A2 U$$58/A1 U$$416/X VGND VGND VPWR VPWR U$$468/A sky130_fd_sc_hd__a22o_1
XU$$478 U$$478/A U$$547/A VGND VGND VPWR VPWR U$$478/X sky130_fd_sc_hd__xor2_1
XU$$489 U$$78/A1 U$$491/A2 U$$80/A1 U$$416/X VGND VGND VPWR VPWR U$$490/A sky130_fd_sc_hd__a22o_1
XFILLER_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_494_ _495_/CLK _494_/D VGND VGND VPWR VPWR _494_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_95_0 dadda_fa_6_95_0/A dadda_fa_6_95_0/B dadda_fa_6_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_96_0/B dadda_fa_7_95_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_30_3 U$$1264/X U$$1397/X U$$1530/X VGND VGND VPWR VPWR dadda_fa_3_31_2/A
+ dadda_fa_3_30_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$990 U$$990/A U$$992/B VGND VGND VPWR VPWR U$$990/X sky130_fd_sc_hd__xor2_1
XFILLER_16_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1140 U$$4291/A1 U$$1200/A2 U$$868/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1141/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1151 U$$1151/A U$$1189/B VGND VGND VPWR VPWR U$$1151/X sky130_fd_sc_hd__xor2_1
XU$$1162 U$$66/A1 U$$1200/A2 U$$68/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1163/A sky130_fd_sc_hd__a22o_1
XU$$1173 U$$1173/A U$$1232/A VGND VGND VPWR VPWR U$$1173/X sky130_fd_sc_hd__xor2_1
XFILLER_188_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1184 U$$88/A1 U$$1218/A2 U$$912/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1185/A sky130_fd_sc_hd__a22o_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1195 U$$1195/A U$$1232/A VGND VGND VPWR VPWR U$$1195/X sky130_fd_sc_hd__xor2_1
X_792__844 VGND VGND VPWR VPWR _792__844/HI U$$4429/B sky130_fd_sc_hd__conb_1
XFILLER_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_833__885 VGND VGND VPWR VPWR _833__885/HI U$$4511/B sky130_fd_sc_hd__conb_1
XFILLER_171_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_82_6 U$$3629/X U$$3762/X U$$3895/X VGND VGND VPWR VPWR dadda_fa_2_83_3/B
+ dadda_fa_2_82_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_75_5 U$$3615/X U$$3748/X U$$3881/X VGND VGND VPWR VPWR dadda_fa_2_76_2/A
+ dadda_fa_2_75_5/A sky130_fd_sc_hd__fa_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_4 U$$4133/X U$$4266/X U$$4399/X VGND VGND VPWR VPWR dadda_fa_2_69_1/CIN
+ dadda_fa_2_68_4/CIN sky130_fd_sc_hd__fa_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_2 dadda_fa_4_38_2/A dadda_fa_4_38_2/B dadda_fa_4_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/CIN dadda_fa_5_38_1/CIN sky130_fd_sc_hd__fa_2
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_3 U$$1330/X U$$1463/X U$$1596/X VGND VGND VPWR VPWR dadda_fa_1_64_6/B
+ dadda_fa_1_63_8/B sky130_fd_sc_hd__fa_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_2 dadda_fa_3_40_2/A dadda_fa_3_40_2/B dadda_fa_3_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/A dadda_fa_4_40_2/B sky130_fd_sc_hd__fa_1
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$370 final_adder.U$$370/A final_adder.U$$370/B VGND VGND VPWR VPWR
+ final_adder.U$$370/X sky130_fd_sc_hd__and2_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _615_/CLK _615_/D VGND VGND VPWR VPWR _615_/Q sky130_fd_sc_hd__dfxtp_4
XU$$220 U$$220/A U$$274/A VGND VGND VPWR VPWR U$$220/X sky130_fd_sc_hd__xor2_1
XFILLER_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_33_1 dadda_fa_3_33_1/A dadda_fa_3_33_1/B dadda_fa_3_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_0/CIN dadda_fa_4_33_2/A sky130_fd_sc_hd__fa_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$231 U$$94/A1 U$$141/X U$$94/B1 U$$142/X VGND VGND VPWR VPWR U$$232/A sky130_fd_sc_hd__a22o_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$242 U$$242/A U$$242/B VGND VGND VPWR VPWR U$$242/X sky130_fd_sc_hd__xor2_1
XFILLER_91_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_10_0 dadda_fa_6_10_0/A dadda_fa_6_10_0/B dadda_fa_6_10_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_11_0/B dadda_fa_7_10_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_26_0 U$$1123/X U$$1256/X U$$1389/X VGND VGND VPWR VPWR dadda_fa_4_27_0/B
+ dadda_fa_4_26_1/CIN sky130_fd_sc_hd__fa_1
XU$$253 U$$938/A1 U$$141/X _607_/Q U$$142/X VGND VGND VPWR VPWR U$$254/A sky130_fd_sc_hd__a22o_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$264 U$$264/A _619_/Q VGND VGND VPWR VPWR U$$264/X sky130_fd_sc_hd__xor2_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$275 _620_/Q VGND VGND VPWR VPWR U$$277/B sky130_fd_sc_hd__inv_1
XFILLER_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_546_ _679_/CLK _546_/D VGND VGND VPWR VPWR _546_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$286 U$$971/A1 U$$278/X U$$12/B1 U$$279/X VGND VGND VPWR VPWR U$$287/A sky130_fd_sc_hd__a22o_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$297 U$$297/A U$$357/B VGND VGND VPWR VPWR U$$297/X sky130_fd_sc_hd__xor2_2
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_477_ _480_/CLK _477_/D VGND VGND VPWR VPWR _477_/Q sky130_fd_sc_hd__dfxtp_1
X_776__828 VGND VGND VPWR VPWR _776__828/HI U$$4397/B sky130_fd_sc_hd__conb_1
XFILLER_158_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_817__869 VGND VGND VPWR VPWR _817__869/HI U$$4479/B sky130_fd_sc_hd__conb_1
XFILLER_139_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3 U$$3/A U$$3/B VGND VGND VPWR VPWR U$$3/X sky130_fd_sc_hd__and2_1
XFILLER_173_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput306 _197_/Q VGND VGND VPWR VPWR o[29] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_5 dadda_fa_2_92_5/A dadda_fa_2_92_5/B dadda_fa_2_92_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_93_2/A dadda_fa_4_92_0/A sky130_fd_sc_hd__fa_2
Xoutput317 _207_/Q VGND VGND VPWR VPWR o[39] sky130_fd_sc_hd__buf_2
XFILLER_154_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput328 _217_/Q VGND VGND VPWR VPWR o[49] sky130_fd_sc_hd__buf_2
XFILLER_5_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput339 _227_/Q VGND VGND VPWR VPWR o[59] sky130_fd_sc_hd__buf_2
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_85_4 dadda_fa_2_85_4/A dadda_fa_2_85_4/B dadda_fa_2_85_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/CIN dadda_fa_3_85_3/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_78_3 dadda_fa_2_78_3/A dadda_fa_2_78_3/B dadda_fa_2_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/B dadda_fa_3_78_3/B sky130_fd_sc_hd__fa_2
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_48_1 dadda_fa_5_48_1/A dadda_fa_5_48_1/B dadda_fa_5_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/B dadda_fa_7_48_0/A sky130_fd_sc_hd__fa_2
XFILLER_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_101_2 U$$3401/X U$$3534/X U$$3667/X VGND VGND VPWR VPWR dadda_fa_3_102_2/B
+ dadda_fa_3_101_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_122_1 input154/X dadda_fa_5_122_1/B dadda_ha_4_122_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_6_123_0/B dadda_fa_7_122_0/A sky130_fd_sc_hd__fa_1
XFILLER_104_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_115_0 dadda_fa_5_115_0/A dadda_fa_5_115_0/B dadda_fa_5_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/A dadda_fa_6_115_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_80_3 U$$2295/X U$$2428/X U$$2561/X VGND VGND VPWR VPWR dadda_fa_2_81_1/CIN
+ dadda_fa_2_80_4/B sky130_fd_sc_hd__fa_1
XFILLER_105_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_73_2 U$$2680/X U$$2813/X U$$2946/X VGND VGND VPWR VPWR dadda_fa_2_74_1/A
+ dadda_fa_2_73_4/A sky130_fd_sc_hd__fa_1
XFILLER_63_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_50_1 dadda_fa_4_50_1/A dadda_fa_4_50_1/B dadda_fa_4_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/B dadda_fa_5_50_1/B sky130_fd_sc_hd__fa_2
Xdadda_fa_1_66_1 U$$2932/X U$$3065/X U$$3198/X VGND VGND VPWR VPWR dadda_fa_2_67_0/CIN
+ dadda_fa_2_66_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_2_100_4 U$$4064/X U$$4197/X VGND VGND VPWR VPWR dadda_fa_3_101_2/CIN dadda_fa_4_100_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_43_0 dadda_fa_4_43_0/A dadda_fa_4_43_0/B dadda_fa_4_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/A dadda_fa_5_43_1/A sky130_fd_sc_hd__fa_1
XFILLER_101_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_0 U$$1588/X U$$1721/X U$$1854/X VGND VGND VPWR VPWR dadda_fa_2_60_0/B
+ dadda_fa_2_59_3/B sky130_fd_sc_hd__fa_2
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _543_/CLK _400_/D VGND VGND VPWR VPWR _400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1909 U$$950/A1 U$$1785/X U$$4514/A1 U$$1786/X VGND VGND VPWR VPWR U$$1910/A sky130_fd_sc_hd__a22o_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_331_ _331_/CLK _331_/D VGND VGND VPWR VPWR _331_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_262_ _267_/CLK _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_193_ _448_/CLK _193_/D VGND VGND VPWR VPWR _193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_95_3 dadda_fa_3_95_3/A dadda_fa_3_95_3/B dadda_fa_3_95_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/B dadda_fa_4_95_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_182_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_88_2 dadda_fa_3_88_2/A dadda_fa_3_88_2/B dadda_fa_3_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/A dadda_fa_4_88_2/B sky130_fd_sc_hd__fa_2
XFILLER_163_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_55_1 U$$516/X U$$649/X VGND VGND VPWR VPWR dadda_fa_1_56_8/A dadda_fa_2_55_0/A
+ sky130_fd_sc_hd__ha_4
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_58_0 dadda_fa_6_58_0/A dadda_fa_6_58_0/B dadda_fa_6_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_59_0/B dadda_fa_7_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4502 U$$4502/A1 U$$4388/X U$$4504/A1 U$$4389/X VGND VGND VPWR VPWR U$$4503/A sky130_fd_sc_hd__a22o_1
XU$$4513 U$$4513/A U$$4513/B VGND VGND VPWR VPWR U$$4513/X sky130_fd_sc_hd__xor2_2
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_61_0 U$$129/X U$$262/X U$$395/X VGND VGND VPWR VPWR dadda_fa_1_62_5/CIN
+ dadda_fa_1_61_7/CIN sky130_fd_sc_hd__fa_2
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$16 U$$16/A1 U$$4/X U$$18/A1 U$$5/X VGND VGND VPWR VPWR U$$17/A sky130_fd_sc_hd__a22o_1
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3801 U$$4486/A1 U$$3703/X U$$787/B1 U$$3704/X VGND VGND VPWR VPWR U$$3802/A sky130_fd_sc_hd__a22o_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3812 U$$3812/A U$$3835/A VGND VGND VPWR VPWR U$$3812/X sky130_fd_sc_hd__xor2_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3823 U$$4508/A1 U$$3703/X _611_/Q U$$3704/X VGND VGND VPWR VPWR U$$3824/A sky130_fd_sc_hd__a22o_1
XU$$27 U$$27/A U$$89/B VGND VGND VPWR VPWR U$$27/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_2 U$$4497/X input148/X dadda_fa_4_117_2/CIN VGND VGND VPWR VPWR dadda_fa_5_118_0/CIN
+ dadda_fa_5_117_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$38 U$$38/A1 U$$4/X U$$40/A1 U$$5/X VGND VGND VPWR VPWR U$$39/A sky130_fd_sc_hd__a22o_1
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3834 U$$3834/A U$$3835/A VGND VGND VPWR VPWR U$$3834/X sky130_fd_sc_hd__xor2_1
XU$$49 U$$49/A U$$9/B VGND VGND VPWR VPWR U$$49/X sky130_fd_sc_hd__xor2_1
XU$$3845 U$$3845/A U$$3893/B VGND VGND VPWR VPWR U$$3845/X sky130_fd_sc_hd__xor2_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3856 U$$979/A1 U$$3840/X U$$22/A1 U$$3841/X VGND VGND VPWR VPWR U$$3857/A sky130_fd_sc_hd__a22o_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3867 U$$3867/A U$$3893/B VGND VGND VPWR VPWR U$$3867/X sky130_fd_sc_hd__xor2_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3878 _569_/Q U$$3970/A2 _570_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3879/A sky130_fd_sc_hd__a22o_1
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3889 U$$3889/A U$$3893/B VGND VGND VPWR VPWR U$$3889/X sky130_fd_sc_hd__xor2_1
XFILLER_166_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_529_ _537_/CLK _529_/D VGND VGND VPWR VPWR _529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_90_2 U$$4044/X U$$4177/X U$$4310/X VGND VGND VPWR VPWR dadda_fa_3_91_1/A
+ dadda_fa_3_90_3/A sky130_fd_sc_hd__fa_1
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_83_1 input238/X dadda_fa_2_83_1/B dadda_fa_2_83_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_84_0/CIN dadda_fa_3_83_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_5_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_60_0 dadda_fa_5_60_0/A dadda_fa_5_60_0/B dadda_fa_5_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/A dadda_fa_6_60_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_76_0 dadda_fa_2_76_0/A dadda_fa_2_76_0/B dadda_fa_2_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/B dadda_fa_3_76_2/B sky130_fd_sc_hd__fa_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_7 U$$3170/X U$$3303/X U$$3436/X VGND VGND VPWR VPWR dadda_fa_2_53_2/CIN
+ dadda_fa_2_52_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_798__850 VGND VGND VPWR VPWR _798__850/HI U$$4441/B sky130_fd_sc_hd__conb_1
XFILLER_24_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_839__891 VGND VGND VPWR VPWR _839__891/HI U$$554/A1 sky130_fd_sc_hd__conb_1
XFILLER_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_98_1 dadda_fa_4_98_1/A dadda_fa_4_98_1/B dadda_fa_4_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/B dadda_fa_5_98_1/B sky130_fd_sc_hd__fa_1
XFILLER_125_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_75_0 dadda_fa_7_75_0/A dadda_fa_7_75_0/B dadda_fa_7_75_0/CIN VGND VGND
+ VPWR VPWR _500_/D _371_/D sky130_fd_sc_hd__fa_1
XFILLER_164_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3108 U$$92/B1 U$$3146/A2 U$$96/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3109/A sky130_fd_sc_hd__a22o_1
XU$$3119 U$$3119/A U$$3129/B VGND VGND VPWR VPWR U$$3119/X sky130_fd_sc_hd__xor2_1
XFILLER_189_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2407 _587_/Q U$$2421/A2 _588_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2408/A sky130_fd_sc_hd__a22o_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2418 U$$2418/A U$$2436/B VGND VGND VPWR VPWR U$$2418/X sky130_fd_sc_hd__xor2_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2429 U$$785/A1 U$$2463/A2 U$$924/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2430/A sky130_fd_sc_hd__a22o_1
XU$$1706 U$$3624/A1 U$$1726/A2 U$$3900/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1707/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1717 U$$1717/A U$$1739/B VGND VGND VPWR VPWR U$$1717/X sky130_fd_sc_hd__xor2_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1728 U$$632/A1 U$$1770/A2 U$$771/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1729/A sky130_fd_sc_hd__a22o_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1739 U$$1739/A U$$1739/B VGND VGND VPWR VPWR U$$1739/X sky130_fd_sc_hd__xor2_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _454_/CLK _314_/D VGND VGND VPWR VPWR _314_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_245_ _503_/CLK _245_/D VGND VGND VPWR VPWR _245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 a[23] VGND VGND VPWR VPWR _639_/D sky130_fd_sc_hd__buf_2
Xinput27 a[33] VGND VGND VPWR VPWR _649_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 a[43] VGND VGND VPWR VPWR _659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_176_ _458_/CLK hold6/X VGND VGND VPWR VPWR _176_/Q sky130_fd_sc_hd__dfxtp_1
Xinput49 a[53] VGND VGND VPWR VPWR _669_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_3_93_0 dadda_fa_3_93_0/A dadda_fa_3_93_0/B dadda_fa_3_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/B dadda_fa_4_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater606 U$$262/B VGND VGND VPWR VPWR U$$242/B sky130_fd_sc_hd__buf_12
XFILLER_81_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater617 _613_/Q VGND VGND VPWR VPWR U$$4514/A1 sky130_fd_sc_hd__buf_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater628 _607_/Q VGND VGND VPWR VPWR U$$940/A1 sky130_fd_sc_hd__buf_12
XU$$4310 U$$4310/A U$$4332/B VGND VGND VPWR VPWR U$$4310/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_55_5 dadda_fa_2_55_5/A dadda_fa_2_55_5/B dadda_fa_2_55_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_2/A dadda_fa_4_55_0/A sky130_fd_sc_hd__fa_2
XFILLER_65_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater639 U$$928/B1 VGND VGND VPWR VPWR U$$4492/A1 sky130_fd_sc_hd__buf_12
XFILLER_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4321 _585_/Q U$$4251/X _586_/Q U$$4252/X VGND VGND VPWR VPWR U$$4322/A sky130_fd_sc_hd__a22o_1
XFILLER_38_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4332 U$$4332/A U$$4332/B VGND VGND VPWR VPWR U$$4332/X sky130_fd_sc_hd__xor2_1
XU$$4343 U$$94/B1 U$$4381/A2 U$$98/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4344/A sky130_fd_sc_hd__a22o_1
XFILLER_19_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4354 U$$4354/A U$$4384/A VGND VGND VPWR VPWR U$$4354/X sky130_fd_sc_hd__xor2_1
XU$$3620 _577_/Q U$$3668/A2 U$$4170/A1 U$$3668/B2 VGND VGND VPWR VPWR U$$3621/A sky130_fd_sc_hd__a22o_1
XU$$4365 U$$4502/A1 U$$4377/A2 U$$4504/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4366/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_4 dadda_fa_2_48_4/A dadda_fa_2_48_4/B dadda_fa_2_48_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/CIN dadda_fa_3_48_3/CIN sky130_fd_sc_hd__fa_1
XU$$3631 U$$3631/A U$$3699/A VGND VGND VPWR VPWR U$$3631/X sky130_fd_sc_hd__xor2_1
XU$$4376 U$$4376/A U$$4384/A VGND VGND VPWR VPWR U$$4376/X sky130_fd_sc_hd__xor2_1
XU$$3642 U$$902/A1 U$$3668/A2 U$$902/B1 U$$3668/B2 VGND VGND VPWR VPWR U$$3643/A sky130_fd_sc_hd__a22o_1
XFILLER_19_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4387 U$$4387/A U$$4387/B VGND VGND VPWR VPWR U$$4387/X sky130_fd_sc_hd__and2_1
XFILLER_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4398 _555_/Q U$$4388/X _556_/Q U$$4389/X VGND VGND VPWR VPWR U$$4399/A sky130_fd_sc_hd__a22o_2
XU$$3653 U$$3653/A U$$3698/A VGND VGND VPWR VPWR U$$3653/X sky130_fd_sc_hd__xor2_1
XU$$3664 U$$4486/A1 U$$3668/A2 _600_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3665/A sky130_fd_sc_hd__a22o_1
XU$$3675 U$$3675/A _669_/Q VGND VGND VPWR VPWR U$$3675/X sky130_fd_sc_hd__xor2_1
XU$$2930 U$$2930/A U$$2996/B VGND VGND VPWR VPWR U$$2930/X sky130_fd_sc_hd__xor2_1
XU$$2941 U$$3900/A1 U$$2975/A2 U$$3489/B1 U$$2975/B2 VGND VGND VPWR VPWR U$$2942/A
+ sky130_fd_sc_hd__a22o_1
XU$$3686 U$$4508/A1 U$$3566/X _611_/Q U$$3567/X VGND VGND VPWR VPWR U$$3687/A sky130_fd_sc_hd__a22o_1
XU$$3697 U$$3697/A U$$3698/A VGND VGND VPWR VPWR U$$3697/X sky130_fd_sc_hd__xor2_1
XU$$2952 U$$2952/A U$$2960/B VGND VGND VPWR VPWR U$$2952/X sky130_fd_sc_hd__xor2_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2963 U$$908/A1 U$$2975/A2 U$$4335/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2964/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2974 U$$2974/A U$$2996/B VGND VGND VPWR VPWR U$$2974/X sky130_fd_sc_hd__xor2_1
XFILLER_34_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2985 U$$4492/A1 U$$2881/X U$$4494/A1 U$$2882/X VGND VGND VPWR VPWR U$$2986/A sky130_fd_sc_hd__a22o_1
XFILLER_179_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2996 U$$2996/A U$$2996/B VGND VGND VPWR VPWR U$$2996/X sky130_fd_sc_hd__xor2_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_44_5 U$$2090/X U$$2223/X VGND VGND VPWR VPWR dadda_fa_2_45_4/A dadda_fa_3_44_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_102_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_50_4 U$$1703/X U$$1836/X U$$1969/X VGND VGND VPWR VPWR dadda_fa_2_51_1/CIN
+ dadda_fa_2_50_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$808 U$$808/A U$$822/A VGND VGND VPWR VPWR U$$808/X sky130_fd_sc_hd__xor2_1
XU$$819 U$$819/A1 U$$689/X U$$819/B1 U$$690/X VGND VGND VPWR VPWR U$$820/A sky130_fd_sc_hd__a22o_1
XFILLER_84_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_43_3 U$$1290/X U$$1423/X U$$1556/X VGND VGND VPWR VPWR dadda_fa_2_44_3/CIN
+ dadda_fa_2_43_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_20_2 dadda_fa_4_20_2/A dadda_fa_4_20_2/B dadda_ha_3_20_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/CIN dadda_fa_5_20_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_13_1 U$$432/X U$$565/X U$$698/X VGND VGND VPWR VPWR dadda_fa_5_14_0/B
+ dadda_fa_5_13_1/B sky130_fd_sc_hd__fa_1
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_58_3 dadda_fa_3_58_3/A dadda_fa_3_58_3/B dadda_fa_3_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/B dadda_fa_4_58_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2204 U$$4122/A1 U$$2270/A2 U$$14/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2205/A sky130_fd_sc_hd__a22o_1
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2215 U$$2215/A U$$2257/B VGND VGND VPWR VPWR U$$2215/X sky130_fd_sc_hd__xor2_1
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2226 U$$3457/B1 U$$2270/A2 U$$4283/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2227/A
+ sky130_fd_sc_hd__a22o_1
XU$$2237 U$$2237/A U$$2257/B VGND VGND VPWR VPWR U$$2237/X sky130_fd_sc_hd__xor2_1
XU$$1503 U$$1503/A _637_/Q VGND VGND VPWR VPWR U$$1503/X sky130_fd_sc_hd__xor2_1
XU$$2248 U$$4303/A1 U$$2270/A2 U$$4442/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2249/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1514 U$$1514/A U$$1614/B VGND VGND VPWR VPWR U$$1514/X sky130_fd_sc_hd__xor2_1
XU$$2259 U$$2259/A U$$2289/B VGND VGND VPWR VPWR U$$2259/X sky130_fd_sc_hd__xor2_1
XFILLER_16_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1525 U$$18/A1 U$$1511/X U$$20/A1 U$$1512/X VGND VGND VPWR VPWR U$$1526/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1536 U$$1536/A U$$1580/B VGND VGND VPWR VPWR U$$1536/X sky130_fd_sc_hd__xor2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1547 U$$3191/A1 U$$1591/A2 U$$3876/B1 U$$1591/B2 VGND VGND VPWR VPWR U$$1548/A
+ sky130_fd_sc_hd__a22o_1
XU$$1558 U$$1558/A U$$1580/B VGND VGND VPWR VPWR U$$1558/X sky130_fd_sc_hd__xor2_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1569 U$$62/A1 U$$1511/X U$$64/A1 U$$1512/X VGND VGND VPWR VPWR U$$1570/A sky130_fd_sc_hd__a22o_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_228_ _499_/CLK _228_/D VGND VGND VPWR VPWR _228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_60_3 dadda_fa_2_60_3/A dadda_fa_2_60_3/B dadda_fa_2_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/B dadda_fa_3_60_3/B sky130_fd_sc_hd__fa_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater403 U$$3703/X VGND VGND VPWR VPWR U$$3783/A2 sky130_fd_sc_hd__buf_12
Xrepeater414 U$$3146/A2 VGND VGND VPWR VPWR U$$3090/A2 sky130_fd_sc_hd__buf_12
Xrepeater425 U$$2470/X VGND VGND VPWR VPWR U$$2574/A2 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_53_2 dadda_fa_2_53_2/A dadda_fa_2_53_2/B dadda_fa_2_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/A dadda_fa_3_53_3/A sky130_fd_sc_hd__fa_1
Xrepeater436 U$$1922/X VGND VGND VPWR VPWR U$$2052/A2 sky130_fd_sc_hd__buf_12
Xrepeater447 U$$1374/X VGND VGND VPWR VPWR U$$1474/A2 sky130_fd_sc_hd__buf_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater458 U$$690/X VGND VGND VPWR VPWR U$$817/B2 sky130_fd_sc_hd__buf_12
XU$$4140 _563_/Q U$$4198/A2 _564_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4141/A sky130_fd_sc_hd__a22o_1
XU$$4151 U$$4151/A U$$4197/B VGND VGND VPWR VPWR U$$4151/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_30_1 dadda_fa_5_30_1/A dadda_fa_5_30_1/B dadda_fa_5_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/B dadda_fa_7_30_0/A sky130_fd_sc_hd__fa_2
Xrepeater469 U$$3678/B2 VGND VGND VPWR VPWR U$$3624/B2 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_46_1 U$$3158/X U$$3224/B input197/X VGND VGND VPWR VPWR dadda_fa_3_47_0/CIN
+ dadda_fa_3_46_2/CIN sky130_fd_sc_hd__fa_1
XU$$4162 _574_/Q U$$4244/A2 U$$4438/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4163/A sky130_fd_sc_hd__a22o_1
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4173 U$$4173/A U$$4197/B VGND VGND VPWR VPWR U$$4173/X sky130_fd_sc_hd__xor2_1
XU$$4184 U$$759/A1 U$$4244/A2 U$$759/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4185/A sky130_fd_sc_hd__a22o_1
XFILLER_66_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_23_0 dadda_fa_5_23_0/A dadda_fa_5_23_0/B dadda_fa_5_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/A dadda_fa_6_23_0/CIN sky130_fd_sc_hd__fa_1
XU$$3450 U$$3450/A U$$3496/B VGND VGND VPWR VPWR U$$3450/X sky130_fd_sc_hd__xor2_1
XU$$4195 U$$4195/A U$$4247/A VGND VGND VPWR VPWR U$$4195/X sky130_fd_sc_hd__xor2_1
XU$$3461 _566_/Q U$$3429/X _567_/Q U$$3430/X VGND VGND VPWR VPWR U$$3462/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_0 U$$1149/X U$$1282/X U$$1415/X VGND VGND VPWR VPWR dadda_fa_3_40_0/B
+ dadda_fa_3_39_2/B sky130_fd_sc_hd__fa_2
XU$$3472 U$$3472/A U$$3496/B VGND VGND VPWR VPWR U$$3472/X sky130_fd_sc_hd__xor2_1
XU$$3483 U$$4442/A1 U$$3429/X _578_/Q U$$3430/X VGND VGND VPWR VPWR U$$3484/A sky130_fd_sc_hd__a22o_1
XFILLER_168_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3494 U$$3494/A U$$3496/B VGND VGND VPWR VPWR U$$3494/X sky130_fd_sc_hd__xor2_1
XU$$2760 U$$979/A1 U$$2796/A2 U$$979/B1 U$$2826/B2 VGND VGND VPWR VPWR U$$2761/A sky130_fd_sc_hd__a22o_1
XU$$2771 U$$2771/A U$$2839/B VGND VGND VPWR VPWR U$$2771/X sky130_fd_sc_hd__xor2_1
XU$$2782 U$$4289/A1 U$$2870/A2 U$$4289/B1 U$$2834/B2 VGND VGND VPWR VPWR U$$2783/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2793 U$$2793/A U$$2797/B VGND VGND VPWR VPWR U$$2793/X sky130_fd_sc_hd__xor2_1
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_68_2 dadda_fa_4_68_2/A dadda_fa_4_68_2/B dadda_fa_4_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/CIN dadda_fa_5_68_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput206 c[54] VGND VGND VPWR VPWR input206/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput217 c[64] VGND VGND VPWR VPWR input217/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput228 c[74] VGND VGND VPWR VPWR input228/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput239 c[84] VGND VGND VPWR VPWR input239/X sky130_fd_sc_hd__buf_2
XFILLER_5_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$700 final_adder.U$$700/A final_adder.U$$700/B VGND VGND VPWR VPWR
+ _246_/D sky130_fd_sc_hd__xor2_1
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$711 final_adder.U$$711/A final_adder.U$$711/B VGND VGND VPWR VPWR
+ _257_/D sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_38_0 dadda_fa_7_38_0/A dadda_fa_7_38_0/B dadda_fa_7_38_0/CIN VGND VGND
+ VPWR VPWR _463_/D _334_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$722 final_adder.U$$722/A final_adder.U$$722/B VGND VGND VPWR VPWR
+ _268_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$733 final_adder.U$$733/A final_adder.U$$733/B VGND VGND VPWR VPWR
+ _279_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$744 final_adder.U$$744/A final_adder.U$$744/B VGND VGND VPWR VPWR
+ _290_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$605 U$$605/A U$$661/B VGND VGND VPWR VPWR U$$605/X sky130_fd_sc_hd__xor2_1
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$616 U$$68/A1 U$$682/A2 U$$68/B1 U$$553/X VGND VGND VPWR VPWR U$$617/A sky130_fd_sc_hd__a22o_1
XFILLER_112_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$627 U$$627/A _625_/Q VGND VGND VPWR VPWR U$$627/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_41_0 U$$89/X U$$222/X U$$355/X VGND VGND VPWR VPWR dadda_fa_2_42_3/B dadda_fa_2_41_5/A
+ sky130_fd_sc_hd__fa_1
XFILLER_186_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$638 U$$90/A1 U$$552/X U$$92/A1 U$$553/X VGND VGND VPWR VPWR U$$639/A sky130_fd_sc_hd__a22o_1
XU$$649 U$$649/A U$$661/B VGND VGND VPWR VPWR U$$649/X sky130_fd_sc_hd__xor2_1
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_70_2 dadda_fa_3_70_2/A dadda_fa_3_70_2/B dadda_fa_3_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/A dadda_fa_4_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_63_1 dadda_fa_3_63_1/A dadda_fa_3_63_1/B dadda_fa_3_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/CIN dadda_fa_4_63_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_40_0 dadda_fa_6_40_0/A dadda_fa_6_40_0/B dadda_fa_6_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_41_0/B dadda_fa_7_40_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_56_0 dadda_fa_3_56_0/A dadda_fa_3_56_0/B dadda_fa_3_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/B dadda_fa_4_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2001 U$$2001/A U$$2021/B VGND VGND VPWR VPWR U$$2001/X sky130_fd_sc_hd__xor2_1
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2012 _595_/Q U$$2036/A2 _596_/Q U$$2036/B2 VGND VGND VPWR VPWR U$$2013/A sky130_fd_sc_hd__a22o_1
XFILLER_63_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_744__796 VGND VGND VPWR VPWR _744__796/HI U$$3020/A1 sky130_fd_sc_hd__conb_1
XU$$2023 U$$2023/A U$$2023/B VGND VGND VPWR VPWR U$$2023/X sky130_fd_sc_hd__xor2_1
XFILLER_35_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2034 _606_/Q U$$2036/A2 _607_/Q U$$2036/B2 VGND VGND VPWR VPWR U$$2035/A sky130_fd_sc_hd__a22o_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2045 U$$2045/A U$$2055/A VGND VGND VPWR VPWR U$$2045/X sky130_fd_sc_hd__xor2_1
XU$$1300 U$$1300/A U$$1342/B VGND VGND VPWR VPWR U$$1300/X sky130_fd_sc_hd__xor2_1
XU$$2056 _646_/Q VGND VGND VPWR VPWR U$$2058/B sky130_fd_sc_hd__inv_1
XU$$1311 U$$76/B1 U$$1367/A2 U$$902/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1312/A sky130_fd_sc_hd__a22o_1
XFILLER_90_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1322 U$$1322/A U$$1369/A VGND VGND VPWR VPWR U$$1322/X sky130_fd_sc_hd__xor2_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2067 U$$12/A1 U$$2117/A2 U$$14/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2068/A sky130_fd_sc_hd__a22o_1
XU$$1333 U$$98/B1 U$$1237/X U$$924/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1334/A sky130_fd_sc_hd__a22o_1
XU$$2078 U$$2078/A U$$2186/B VGND VGND VPWR VPWR U$$2078/X sky130_fd_sc_hd__xor2_1
XU$$2089 U$$3457/B1 U$$2117/A2 U$$4283/A1 U$$2117/B2 VGND VGND VPWR VPWR U$$2090/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1344 U$$1344/A U$$1369/A VGND VGND VPWR VPWR U$$1344/X sky130_fd_sc_hd__xor2_1
XU$$1355 U$$944/A1 U$$1367/A2 U$$946/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1356/A sky130_fd_sc_hd__a22o_1
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1366 U$$1366/A U$$1369/A VGND VGND VPWR VPWR U$$1366/X sky130_fd_sc_hd__xor2_1
XU$$1377 U$$1377/A U$$1479/B VGND VGND VPWR VPWR U$$1377/X sky130_fd_sc_hd__xor2_1
XFILLER_188_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1388 U$$18/A1 U$$1474/A2 U$$20/A1 U$$1466/B2 VGND VGND VPWR VPWR U$$1389/A sky130_fd_sc_hd__a22o_1
XU$$1399 U$$1399/A U$$1479/B VGND VGND VPWR VPWR U$$1399/X sky130_fd_sc_hd__xor2_1
XFILLER_148_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_113_0 dadda_fa_7_113_0/A dadda_fa_7_113_0/B dadda_fa_7_113_0/CIN VGND
+ VGND VPWR VPWR _538_/D _409_/D sky130_fd_sc_hd__fa_2
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_78_1 dadda_fa_5_78_1/A dadda_fa_5_78_1/B dadda_fa_5_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/B dadda_fa_7_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_135_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$40 _464_/Q _336_/Q VGND VGND VPWR VPWR final_adder.U$$535/B1 final_adder.U$$662/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$51 _475_/Q _347_/Q VGND VGND VPWR VPWR final_adder.U$$179/B1 final_adder.U$$673/A
+ sky130_fd_sc_hd__ha_1
XU$$3280 U$$3280/A _663_/Q VGND VGND VPWR VPWR U$$3280/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$62 _486_/Q _358_/Q VGND VGND VPWR VPWR final_adder.U$$557/B1 final_adder.U$$684/A
+ sky130_fd_sc_hd__ha_1
XU$$3291 _665_/Q U$$3291/B VGND VGND VPWR VPWR U$$3291/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$73 _497_/Q _369_/Q VGND VGND VPWR VPWR final_adder.U$$201/B1 final_adder.U$$695/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$84 _508_/Q _380_/Q VGND VGND VPWR VPWR final_adder.U$$579/B1 final_adder.U$$706/A
+ sky130_fd_sc_hd__ha_1
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$95 _519_/Q _391_/Q VGND VGND VPWR VPWR final_adder.U$$223/B1 final_adder.U$$717/A
+ sky130_fd_sc_hd__ha_1
XU$$2590 _610_/Q U$$2470/X _611_/Q U$$2471/X VGND VGND VPWR VPWR U$$2591/A sky130_fd_sc_hd__a22o_1
XFILLER_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_693__913 VGND VGND VPWR VPWR _693__913/HI _693__913/LO sky130_fd_sc_hd__conb_1
XFILLER_22_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_80_1 dadda_fa_4_80_1/A dadda_fa_4_80_1/B dadda_fa_4_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/B dadda_fa_5_80_1/B sky130_fd_sc_hd__fa_1
XFILLER_135_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_73_0 dadda_fa_4_73_0/A dadda_fa_4_73_0/B dadda_fa_4_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/A dadda_fa_5_73_1/A sky130_fd_sc_hd__fa_1
XFILLER_122_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_89_0 U$$1780/Y U$$1914/X U$$2047/X VGND VGND VPWR VPWR dadda_fa_2_90_3/CIN
+ dadda_fa_2_89_5/A sky130_fd_sc_hd__fa_2
XFILLER_66_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$541 final_adder.U$$668/A final_adder.U$$668/B final_adder.U$$541/B1
+ VGND VGND VPWR VPWR final_adder.U$$669/B sky130_fd_sc_hd__a21o_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_631_ _646_/CLK _631_/D VGND VGND VPWR VPWR _631_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$563 final_adder.U$$690/A final_adder.U$$690/B final_adder.U$$563/B1
+ VGND VGND VPWR VPWR final_adder.U$$691/B sky130_fd_sc_hd__a21o_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$402 U$$539/A1 U$$278/X U$$952/A1 U$$279/X VGND VGND VPWR VPWR U$$403/A sky130_fd_sc_hd__a22o_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$413 _623_/Q VGND VGND VPWR VPWR U$$413/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$585 final_adder.U$$712/A final_adder.U$$712/B final_adder.U$$585/B1
+ VGND VGND VPWR VPWR final_adder.U$$713/B sky130_fd_sc_hd__a21o_1
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$424 U$$424/A U$$530/B VGND VGND VPWR VPWR U$$424/X sky130_fd_sc_hd__xor2_1
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$435 _560_/Q U$$491/A2 U$$26/A1 U$$416/X VGND VGND VPWR VPWR U$$436/A sky130_fd_sc_hd__a22o_1
XFILLER_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_562_ _637_/CLK _562_/D VGND VGND VPWR VPWR _562_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$446 U$$446/A U$$530/B VGND VGND VPWR VPWR U$$446/X sky130_fd_sc_hd__xor2_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$457 U$$46/A1 U$$491/A2 _572_/Q U$$416/X VGND VGND VPWR VPWR U$$458/A sky130_fd_sc_hd__a22o_1
XU$$468 U$$468/A U$$530/B VGND VGND VPWR VPWR U$$468/X sky130_fd_sc_hd__xor2_1
XFILLER_32_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$479 U$$68/A1 U$$491/A2 U$$68/B1 U$$416/X VGND VGND VPWR VPWR U$$480/A sky130_fd_sc_hd__a22o_1
X_493_ _496_/CLK _493_/D VGND VGND VPWR VPWR _493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_88_0 dadda_fa_6_88_0/A dadda_fa_6_88_0/B dadda_fa_6_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_89_0/B dadda_fa_7_88_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_78_0 _704__924/HI U$$1094/X VGND VGND VPWR VPWR dadda_fa_2_79_0/A dadda_fa_2_78_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$980 U$$980/A U$$980/B VGND VGND VPWR VPWR U$$980/X sky130_fd_sc_hd__xor2_2
XU$$1130 U$$34/A1 U$$1100/X U$$36/A1 U$$1101/X VGND VGND VPWR VPWR U$$1131/A sky130_fd_sc_hd__a22o_1
XU$$991 U$$32/A1 U$$999/A2 U$$34/A1 U$$999/B2 VGND VGND VPWR VPWR U$$992/A sky130_fd_sc_hd__a22o_1
XU$$1141 U$$1141/A U$$1167/B VGND VGND VPWR VPWR U$$1141/X sky130_fd_sc_hd__xor2_1
XU$$1152 U$$56/A1 U$$1100/X U$$58/A1 U$$1101/X VGND VGND VPWR VPWR U$$1153/A sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1163 U$$1163/A U$$1167/B VGND VGND VPWR VPWR U$$1163/X sky130_fd_sc_hd__xor2_1
XFILLER_176_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1174 U$$76/B1 U$$1218/A2 U$$902/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1175/A sky130_fd_sc_hd__a22o_1
XU$$1185 U$$1185/A U$$1232/A VGND VGND VPWR VPWR U$$1185/X sky130_fd_sc_hd__xor2_1
XU$$1196 U$$98/B1 U$$1218/A2 U$$924/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1197/A sky130_fd_sc_hd__a22o_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_90_0 dadda_fa_5_90_0/A dadda_fa_5_90_0/B dadda_fa_5_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/A dadda_fa_6_90_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_75_6 U$$4014/X U$$4147/X U$$4280/X VGND VGND VPWR VPWR dadda_fa_2_76_2/B
+ dadda_fa_2_75_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_68_5 input221/X dadda_fa_1_68_5/B dadda_fa_1_68_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_69_2/A dadda_fa_2_68_5/A sky130_fd_sc_hd__fa_2
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_120_0 dadda_fa_6_120_0/A dadda_fa_6_120_0/B dadda_fa_6_120_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_121_0/B dadda_fa_7_120_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_7_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_4 U$$1729/X U$$1862/X U$$1995/X VGND VGND VPWR VPWR dadda_fa_1_64_6/CIN
+ dadda_fa_1_63_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_40_3 dadda_fa_3_40_3/A dadda_fa_3_40_3/B dadda_fa_3_40_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/B dadda_fa_4_40_2/CIN sky130_fd_sc_hd__fa_2
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$360 final_adder.U$$360/A final_adder.U$$360/B VGND VGND VPWR VPWR
+ final_adder.U$$372/B sky130_fd_sc_hd__and2_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$371 final_adder.U$$370/A final_adder.U$$357/X final_adder.U$$359/X
+ VGND VGND VPWR VPWR final_adder.U$$371/X sky130_fd_sc_hd__a21o_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$210 U$$210/A U$$242/B VGND VGND VPWR VPWR U$$210/X sky130_fd_sc_hd__xor2_1
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$221 U$$84/A1 U$$141/X U$$86/A1 U$$142/X VGND VGND VPWR VPWR U$$222/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_33_2 dadda_fa_3_33_2/A dadda_fa_3_33_2/B dadda_fa_3_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/A dadda_fa_4_33_2/B sky130_fd_sc_hd__fa_2
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_614_ _614_/CLK _614_/D VGND VGND VPWR VPWR _614_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$393 final_adder.U$$356/B final_adder.U$$654/B final_adder.U$$329/X
+ VGND VGND VPWR VPWR final_adder.U$$662/B sky130_fd_sc_hd__a21o_2
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$232 U$$232/A U$$274/A VGND VGND VPWR VPWR U$$232/X sky130_fd_sc_hd__xor2_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$243 U$$928/A1 U$$141/X U$$928/B1 U$$142/X VGND VGND VPWR VPWR U$$244/A sky130_fd_sc_hd__a22o_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$254 U$$254/A U$$262/B VGND VGND VPWR VPWR U$$254/X sky130_fd_sc_hd__xor2_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$265 U$$539/A1 U$$141/X U$$952/A1 U$$142/X VGND VGND VPWR VPWR U$$266/A sky130_fd_sc_hd__a22o_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_26_1 U$$1522/X U$$1655/X U$$1788/X VGND VGND VPWR VPWR dadda_fa_4_27_0/CIN
+ dadda_fa_4_26_2/A sky130_fd_sc_hd__fa_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_545_ _598_/CLK _545_/D VGND VGND VPWR VPWR _545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$276 _621_/Q VGND VGND VPWR VPWR U$$276/Y sky130_fd_sc_hd__inv_1
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$287 U$$287/A U$$357/B VGND VGND VPWR VPWR U$$287/X sky130_fd_sc_hd__xor2_1
XFILLER_72_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$298 U$$983/A1 U$$278/X _561_/Q U$$279/X VGND VGND VPWR VPWR U$$299/A sky130_fd_sc_hd__a22o_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_19_0 U$$45/X U$$178/X U$$311/X VGND VGND VPWR VPWR dadda_fa_4_20_0/CIN
+ dadda_fa_4_19_2/A sky130_fd_sc_hd__fa_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ _476_/CLK _476_/D VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4 U$$2/Y U$$1/A U$$4/A3 U$$3/X U$$0/Y VGND VGND VPWR VPWR U$$4/X sky130_fd_sc_hd__a32o_4
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput307 _170_/Q VGND VGND VPWR VPWR o[2] sky130_fd_sc_hd__buf_2
Xoutput318 _171_/Q VGND VGND VPWR VPWR o[3] sky130_fd_sc_hd__buf_2
Xoutput329 _172_/Q VGND VGND VPWR VPWR o[4] sky130_fd_sc_hd__buf_2
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_85_5 dadda_fa_2_85_5/A dadda_fa_2_85_5/B dadda_fa_2_85_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_2/A dadda_fa_4_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_78_4 dadda_fa_2_78_4/A dadda_fa_2_78_4/B dadda_fa_2_78_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/CIN dadda_fa_3_78_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_141_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_101_3 U$$3800/X U$$3933/X U$$4066/X VGND VGND VPWR VPWR dadda_fa_3_102_2/CIN
+ dadda_fa_4_101_0/A sky130_fd_sc_hd__fa_1
XFILLER_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_800__852 VGND VGND VPWR VPWR _800__852/HI U$$4445/B sky130_fd_sc_hd__conb_1
XFILLER_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_115_1 dadda_fa_5_115_1/A dadda_fa_5_115_1/B dadda_fa_5_115_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/B dadda_fa_7_115_0/A sky130_fd_sc_hd__fa_1
XFILLER_176_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_108_0 dadda_fa_5_108_0/A dadda_fa_5_108_0/B dadda_fa_5_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/A dadda_fa_6_108_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_80_4 U$$2694/X U$$2827/X U$$2960/X VGND VGND VPWR VPWR dadda_fa_2_81_2/A
+ dadda_fa_2_80_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_63_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_73_3 U$$3079/X U$$3212/X U$$3345/X VGND VGND VPWR VPWR dadda_fa_2_74_1/B
+ dadda_fa_2_73_4/B sky130_fd_sc_hd__fa_1
XFILLER_59_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_50_2 dadda_fa_4_50_2/A dadda_fa_4_50_2/B dadda_fa_4_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/CIN dadda_fa_5_50_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_66_2 U$$3331/X U$$3464/X U$$3597/X VGND VGND VPWR VPWR dadda_fa_2_67_1/A
+ dadda_fa_2_66_4/A sky130_fd_sc_hd__fa_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_43_1 dadda_fa_4_43_1/A dadda_fa_4_43_1/B dadda_fa_4_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/B dadda_fa_5_43_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_59_1 U$$1987/X U$$2120/X U$$2253/X VGND VGND VPWR VPWR dadda_fa_2_60_0/CIN
+ dadda_fa_2_59_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_132_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_20_0 dadda_fa_7_20_0/A dadda_fa_7_20_0/B dadda_fa_7_20_0/CIN VGND VGND
+ VPWR VPWR _445_/D _316_/D sky130_fd_sc_hd__fa_2
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_36_0 dadda_fa_4_36_0/A dadda_fa_4_36_0/B dadda_fa_4_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/A dadda_fa_5_36_1/A sky130_fd_sc_hd__fa_1
XFILLER_55_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_330_ _333_/CLK _330_/D VGND VGND VPWR VPWR _330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _280_/CLK _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_192_ _448_/CLK _192_/D VGND VGND VPWR VPWR _192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_88_3 dadda_fa_3_88_3/A dadda_fa_3_88_3/B dadda_fa_3_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/B dadda_fa_4_88_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_163_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4503 U$$4503/A U$$4503/B VGND VGND VPWR VPWR U$$4503/X sky130_fd_sc_hd__xor2_2
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4514 U$$4514/A1 U$$4388/X U$$952/B1 U$$4389/X VGND VGND VPWR VPWR U$$4515/A sky130_fd_sc_hd__a22o_1
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_61_1 U$$528/X U$$661/X U$$794/X VGND VGND VPWR VPWR dadda_fa_1_62_6/A
+ dadda_fa_1_61_8/A sky130_fd_sc_hd__fa_1
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$17 U$$17/A U$$9/B VGND VGND VPWR VPWR U$$17/X sky130_fd_sc_hd__xor2_1
XU$$3802 U$$3802/A U$$3835/A VGND VGND VPWR VPWR U$$3802/X sky130_fd_sc_hd__xor2_1
XU$$28 U$$28/A1 U$$4/X U$$28/B1 U$$5/X VGND VGND VPWR VPWR U$$29/A sky130_fd_sc_hd__a22o_1
XU$$3813 _605_/Q U$$3703/X U$$4500/A1 U$$3704/X VGND VGND VPWR VPWR U$$3814/A sky130_fd_sc_hd__a22o_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3824 U$$3824/A U$$3835/A VGND VGND VPWR VPWR U$$3824/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_54_0 U$$115/X U$$248/X U$$381/X VGND VGND VPWR VPWR dadda_fa_1_55_8/A
+ dadda_fa_1_54_8/CIN sky130_fd_sc_hd__fa_2
XFILLER_58_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$39 U$$39/A U$$3/A VGND VGND VPWR VPWR U$$39/X sky130_fd_sc_hd__xor2_1
XU$$3835 U$$3835/A VGND VGND VPWR VPWR U$$3835/Y sky130_fd_sc_hd__inv_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3846 _553_/Q U$$3912/A2 U$$4122/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3847/A sky130_fd_sc_hd__a22o_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$190 final_adder.U$$685/A final_adder.U$$684/A VGND VGND VPWR VPWR
+ final_adder.U$$286/A sky130_fd_sc_hd__and2_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3857 U$$3857/A U$$3929/B VGND VGND VPWR VPWR U$$3857/X sky130_fd_sc_hd__xor2_1
XFILLER_46_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3868 _564_/Q U$$3840/X _565_/Q U$$3841/X VGND VGND VPWR VPWR U$$3869/A sky130_fd_sc_hd__a22o_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3879 U$$3879/A U$$3969/B VGND VGND VPWR VPWR U$$3879/X sky130_fd_sc_hd__xor2_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_528_ _543_/CLK _528_/D VGND VGND VPWR VPWR _528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_459_ _463_/CLK _459_/D VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_90_3 U$$4443/X input246/X dadda_fa_2_90_3/CIN VGND VGND VPWR VPWR dadda_fa_3_91_1/B
+ dadda_fa_3_90_3/B sky130_fd_sc_hd__fa_2
XFILLER_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_83_2 dadda_fa_2_83_2/A dadda_fa_2_83_2/B dadda_fa_2_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/A dadda_fa_3_83_3/A sky130_fd_sc_hd__fa_1
XFILLER_126_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_60_1 dadda_fa_5_60_1/A dadda_fa_5_60_1/B dadda_fa_5_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/B dadda_fa_7_60_0/A sky130_fd_sc_hd__fa_1
XFILLER_130_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_1 dadda_fa_2_76_1/A dadda_fa_2_76_1/B dadda_fa_2_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/CIN dadda_fa_3_76_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_53_0 dadda_fa_5_53_0/A dadda_fa_5_53_0/B dadda_fa_5_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/A dadda_fa_6_53_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_69_0 dadda_fa_2_69_0/A dadda_fa_2_69_0/B dadda_fa_2_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/B dadda_fa_3_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_52_8 U$$3569/X U$$3698/A input204/X VGND VGND VPWR VPWR dadda_fa_2_53_3/A
+ dadda_fa_3_52_0/A sky130_fd_sc_hd__fa_2
XFILLER_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_98_2 dadda_fa_4_98_2/A dadda_fa_4_98_2/B dadda_fa_4_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/CIN dadda_fa_5_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_30_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_68_0 dadda_fa_7_68_0/A dadda_fa_7_68_0/B dadda_fa_7_68_0/CIN VGND VGND
+ VPWR VPWR _493_/D _364_/D sky130_fd_sc_hd__fa_2
XFILLER_160_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_0 U$$2144/X U$$2277/X U$$2410/X VGND VGND VPWR VPWR dadda_fa_2_72_0/B
+ dadda_fa_2_71_3/B sky130_fd_sc_hd__fa_2
XFILLER_87_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3109 U$$3109/A U$$3109/B VGND VGND VPWR VPWR U$$3109/X sky130_fd_sc_hd__xor2_1
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2408 U$$2408/A U$$2436/B VGND VGND VPWR VPWR U$$2408/X sky130_fd_sc_hd__xor2_1
XFILLER_43_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2419 U$$912/A1 U$$2463/A2 U$$914/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2420/A sky130_fd_sc_hd__a22o_1
XFILLER_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1707 U$$1707/A U$$1739/B VGND VGND VPWR VPWR U$$1707/X sky130_fd_sc_hd__xor2_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1718 U$$74/A1 U$$1726/A2 U$$2953/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1719/A sky130_fd_sc_hd__a22o_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1729 U$$1729/A U$$1781/A VGND VGND VPWR VPWR U$$1729/X sky130_fd_sc_hd__xor2_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _463_/CLK _313_/D VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_244_ _503_/CLK _244_/D VGND VGND VPWR VPWR _244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 a[24] VGND VGND VPWR VPWR _640_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_161_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput28 a[34] VGND VGND VPWR VPWR _650_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput39 a[44] VGND VGND VPWR VPWR _660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_175_ _333_/CLK hold3/X VGND VGND VPWR VPWR _175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_93_1 dadda_fa_3_93_1/A dadda_fa_3_93_1/B dadda_fa_3_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/CIN dadda_fa_4_93_2/A sky130_fd_sc_hd__fa_2
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_70_0 dadda_fa_6_70_0/A dadda_fa_6_70_0/B dadda_fa_6_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_71_0/B dadda_fa_7_70_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_86_0 dadda_fa_3_86_0/A dadda_fa_3_86_0/B dadda_fa_3_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/B dadda_fa_4_86_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_124_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater607 U$$262/B VGND VGND VPWR VPWR U$$274/A sky130_fd_sc_hd__buf_12
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4300 U$$4300/A U$$4384/A VGND VGND VPWR VPWR U$$4300/X sky130_fd_sc_hd__xor2_1
Xrepeater618 U$$950/A1 VGND VGND VPWR VPWR U$$539/A1 sky130_fd_sc_hd__buf_12
Xrepeater629 _607_/Q VGND VGND VPWR VPWR U$$4502/A1 sky130_fd_sc_hd__buf_12
XU$$4311 _580_/Q U$$4377/A2 _581_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4312/A sky130_fd_sc_hd__a22o_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4322 U$$4322/A U$$4332/B VGND VGND VPWR VPWR U$$4322/X sky130_fd_sc_hd__xor2_1
XU$$4333 U$$771/A1 U$$4381/A2 _592_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4334/A sky130_fd_sc_hd__a22o_1
XFILLER_120_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4344 U$$4344/A _679_/Q VGND VGND VPWR VPWR U$$4344/X sky130_fd_sc_hd__xor2_1
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3610 U$$4156/B1 U$$3668/A2 _573_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3611/A sky130_fd_sc_hd__a22o_1
XU$$4355 U$$4492/A1 U$$4381/A2 U$$4494/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4356/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3621 U$$3621/A U$$3699/A VGND VGND VPWR VPWR U$$3621/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_0 U$$3961/X U$$4094/X U$$4227/X VGND VGND VPWR VPWR dadda_fa_5_116_0/A
+ dadda_fa_5_115_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_48_5 dadda_fa_2_48_5/A dadda_fa_2_48_5/B dadda_fa_2_48_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_2/A dadda_fa_4_48_0/A sky130_fd_sc_hd__fa_1
XU$$4366 U$$4366/A U$$4384/A VGND VGND VPWR VPWR U$$4366/X sky130_fd_sc_hd__xor2_1
XU$$3632 _583_/Q U$$3668/A2 _584_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3633/A sky130_fd_sc_hd__a22o_1
XU$$4377 _613_/Q U$$4377/A2 U$$4379/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4378/A sky130_fd_sc_hd__a22o_1
XU$$3643 U$$3643/A U$$3699/A VGND VGND VPWR VPWR U$$3643/X sky130_fd_sc_hd__xor2_1
XU$$4388 U$$4386/Y U$$4388/A2 U$$4384/A U$$4387/X U$$4384/Y VGND VGND VPWR VPWR U$$4388/X
+ sky130_fd_sc_hd__a32o_1
XU$$4399 U$$4399/A U$$4399/B VGND VGND VPWR VPWR U$$4399/X sky130_fd_sc_hd__xor2_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3654 _594_/Q U$$3668/A2 _595_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3655/A sky130_fd_sc_hd__a22o_1
XU$$2920 U$$2920/A U$$2960/B VGND VGND VPWR VPWR U$$2920/X sky130_fd_sc_hd__xor2_1
XU$$3665 U$$3665/A U$$3699/A VGND VGND VPWR VPWR U$$3665/X sky130_fd_sc_hd__xor2_1
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2931 U$$54/A1 U$$3009/A2 U$$56/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2932/A sky130_fd_sc_hd__a22o_1
XFILLER_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3676 _605_/Q U$$3566/X U$$4500/A1 U$$3567/X VGND VGND VPWR VPWR U$$3677/A sky130_fd_sc_hd__a22o_1
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2942 U$$2942/A U$$2960/B VGND VGND VPWR VPWR U$$2942/X sky130_fd_sc_hd__xor2_1
XFILLER_18_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3687 U$$3687/A U$$3698/A VGND VGND VPWR VPWR U$$3687/X sky130_fd_sc_hd__xor2_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2953 U$$2953/A1 U$$2975/A2 U$$76/B1 U$$2975/B2 VGND VGND VPWR VPWR U$$2954/A sky130_fd_sc_hd__a22o_1
XU$$3698 U$$3698/A VGND VGND VPWR VPWR U$$3698/Y sky130_fd_sc_hd__inv_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2964 U$$2964/A _659_/Q VGND VGND VPWR VPWR U$$2964/X sky130_fd_sc_hd__xor2_1
XU$$2975 _597_/Q U$$2975/A2 U$$4484/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2976/A sky130_fd_sc_hd__a22o_1
XU$$2986 U$$2986/A _659_/Q VGND VGND VPWR VPWR U$$2986/X sky130_fd_sc_hd__xor2_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2997 _608_/Q U$$2881/X U$$4506/A1 U$$2882/X VGND VGND VPWR VPWR U$$2998/A sky130_fd_sc_hd__a22o_1
XFILLER_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_50_5 U$$2102/X U$$2235/X U$$2368/X VGND VGND VPWR VPWR dadda_fa_2_51_2/A
+ dadda_fa_2_50_5/A sky130_fd_sc_hd__fa_2
XU$$809 U$$946/A1 U$$817/A2 U$$948/A1 U$$817/B2 VGND VGND VPWR VPWR U$$810/A sky130_fd_sc_hd__a22o_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2205 U$$2205/A U$$2257/B VGND VGND VPWR VPWR U$$2205/X sky130_fd_sc_hd__xor2_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2216 U$$983/A1 U$$2270/A2 U$$26/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2217/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2227 U$$2227/A U$$2257/B VGND VGND VPWR VPWR U$$2227/X sky130_fd_sc_hd__xor2_1
XU$$2238 U$$4291/B1 U$$2270/A2 U$$48/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2239/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2249 U$$2249/A U$$2257/B VGND VGND VPWR VPWR U$$2249/X sky130_fd_sc_hd__xor2_1
XU$$1504 _615_/Q U$$1374/X U$$1504/B1 U$$1375/X VGND VGND VPWR VPWR U$$1505/A sky130_fd_sc_hd__a22o_1
XFILLER_90_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1515 U$$8/A1 U$$1511/X U$$8/B1 U$$1512/X VGND VGND VPWR VPWR U$$1516/A sky130_fd_sc_hd__a22o_1
XFILLER_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1526 U$$1526/A U$$1614/B VGND VGND VPWR VPWR U$$1526/X sky130_fd_sc_hd__xor2_1
XFILLER_188_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1537 U$$30/A1 U$$1591/A2 U$$30/B1 U$$1591/B2 VGND VGND VPWR VPWR U$$1538/A sky130_fd_sc_hd__a22o_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1548 U$$1548/A U$$1580/B VGND VGND VPWR VPWR U$$1548/X sky130_fd_sc_hd__xor2_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1559 U$$2790/B1 U$$1605/A2 U$$876/A1 U$$1605/B2 VGND VGND VPWR VPWR U$$1560/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ _474_/CLK _227_/D VGND VGND VPWR VPWR _227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_749__801 VGND VGND VPWR VPWR _749__801/HI U$$3422/B1 sky130_fd_sc_hd__conb_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_60_4 dadda_fa_2_60_4/A dadda_fa_2_60_4/B dadda_fa_2_60_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/CIN dadda_fa_3_60_3/CIN sky130_fd_sc_hd__fa_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater404 U$$3703/X VGND VGND VPWR VPWR U$$3795/A2 sky130_fd_sc_hd__buf_12
XFILLER_111_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater415 U$$3018/X VGND VGND VPWR VPWR U$$3146/A2 sky130_fd_sc_hd__buf_12
Xrepeater426 U$$2463/A2 VGND VGND VPWR VPWR U$$2421/A2 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_53_3 dadda_fa_2_53_3/A dadda_fa_2_53_3/B dadda_fa_2_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/B dadda_fa_3_53_3/B sky130_fd_sc_hd__fa_2
Xrepeater437 U$$1897/A2 VGND VGND VPWR VPWR U$$1903/A2 sky130_fd_sc_hd__buf_12
Xrepeater448 U$$1237/X VGND VGND VPWR VPWR U$$1341/A2 sky130_fd_sc_hd__buf_12
XU$$4130 _558_/Q U$$4244/A2 _559_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4131/A sky130_fd_sc_hd__a22o_1
Xrepeater459 U$$4381/B2 VGND VGND VPWR VPWR U$$4377/B2 sky130_fd_sc_hd__buf_12
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4141 U$$4141/A U$$4247/A VGND VGND VPWR VPWR U$$4141/X sky130_fd_sc_hd__xor2_1
XU$$4152 U$$4289/A1 U$$4114/X U$$4289/B1 U$$4198/B2 VGND VGND VPWR VPWR U$$4153/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4163 U$$4163/A _677_/Q VGND VGND VPWR VPWR U$$4163/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_2 dadda_fa_2_46_2/A dadda_fa_2_46_2/B dadda_fa_2_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/A dadda_fa_3_46_3/A sky130_fd_sc_hd__fa_2
XFILLER_66_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4174 _580_/Q U$$4198/A2 _581_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4175/A sky130_fd_sc_hd__a22o_1
XU$$3440 U$$3440/A U$$3496/B VGND VGND VPWR VPWR U$$3440/X sky130_fd_sc_hd__xor2_1
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4185 U$$4185/A U$$4246/A VGND VGND VPWR VPWR U$$4185/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_23_1 dadda_fa_5_23_1/A dadda_fa_5_23_1/B dadda_fa_5_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/B dadda_fa_7_23_0/A sky130_fd_sc_hd__fa_2
XFILLER_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4196 U$$771/A1 U$$4114/X U$$4335/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4197/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_1 U$$1548/X U$$1681/X U$$1814/X VGND VGND VPWR VPWR dadda_fa_3_40_0/CIN
+ dadda_fa_3_39_2/CIN sky130_fd_sc_hd__fa_2
XU$$3451 U$$4273/A1 U$$3525/A2 U$$28/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3452/A sky130_fd_sc_hd__a22o_1
XU$$3462 U$$3462/A _667_/Q VGND VGND VPWR VPWR U$$3462/X sky130_fd_sc_hd__xor2_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3473 U$$4156/B1 U$$3525/A2 _573_/Q U$$3525/B2 VGND VGND VPWR VPWR U$$3474/A sky130_fd_sc_hd__a22o_1
XFILLER_92_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3484 U$$3484/A U$$3561/A VGND VGND VPWR VPWR U$$3484/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_16_0 dadda_fa_5_16_0/A dadda_fa_5_16_0/B dadda_fa_5_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/A dadda_fa_6_16_0/CIN sky130_fd_sc_hd__fa_1
XU$$2750 U$$969/A1 U$$2796/A2 U$$971/A1 U$$2745/X VGND VGND VPWR VPWR U$$2751/A sky130_fd_sc_hd__a22o_1
XFILLER_179_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3495 U$$892/A1 U$$3525/A2 U$$892/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3496/A sky130_fd_sc_hd__a22o_1
XU$$2761 U$$2761/A U$$2797/B VGND VGND VPWR VPWR U$$2761/X sky130_fd_sc_hd__xor2_1
XU$$2772 _564_/Q U$$2796/A2 _565_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2773/A sky130_fd_sc_hd__a22o_1
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2783 U$$2783/A U$$2839/B VGND VGND VPWR VPWR U$$2783/X sky130_fd_sc_hd__xor2_1
XFILLER_179_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2794 U$$54/A1 U$$2796/A2 U$$56/A1 U$$2745/X VGND VGND VPWR VPWR U$$2795/A sky130_fd_sc_hd__a22o_1
XFILLER_21_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput207 c[55] VGND VGND VPWR VPWR input207/X sky130_fd_sc_hd__buf_2
Xinput218 c[65] VGND VGND VPWR VPWR input218/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput229 c[75] VGND VGND VPWR VPWR input229/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$701 final_adder.U$$701/A final_adder.U$$701/B VGND VGND VPWR VPWR
+ _247_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$712 final_adder.U$$712/A final_adder.U$$712/B VGND VGND VPWR VPWR
+ _258_/D sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$723 final_adder.U$$723/A final_adder.U$$723/B VGND VGND VPWR VPWR
+ _269_/D sky130_fd_sc_hd__xor2_1
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$734 final_adder.U$$734/A final_adder.U$$734/B VGND VGND VPWR VPWR
+ _280_/D sky130_fd_sc_hd__xor2_1
XFILLER_151_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$745 final_adder.U$$745/A final_adder.U$$745/B VGND VGND VPWR VPWR
+ _291_/D sky130_fd_sc_hd__xor2_2
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$606 U$$58/A1 U$$682/A2 U$$60/A1 U$$553/X VGND VGND VPWR VPWR U$$607/A sky130_fd_sc_hd__a22o_1
XU$$617 U$$617/A U$$661/B VGND VGND VPWR VPWR U$$617/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_41_1 U$$488/X U$$621/X U$$754/X VGND VGND VPWR VPWR dadda_fa_2_42_3/CIN
+ dadda_fa_2_41_5/B sky130_fd_sc_hd__fa_1
XU$$628 U$$902/A1 U$$682/A2 U$$902/B1 U$$553/X VGND VGND VPWR VPWR U$$629/A sky130_fd_sc_hd__a22o_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$639 U$$639/A _625_/Q VGND VGND VPWR VPWR U$$639/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_3 dadda_fa_3_70_3/A dadda_fa_3_70_3/B dadda_fa_3_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/B dadda_fa_4_70_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_63_2 dadda_fa_3_63_2/A dadda_fa_3_63_2/B dadda_fa_3_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/A dadda_fa_4_63_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_56_1 dadda_fa_3_56_1/A dadda_fa_3_56_1/B dadda_fa_3_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/CIN dadda_fa_4_56_2/A sky130_fd_sc_hd__fa_1
XFILLER_94_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_43_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_33_0 dadda_fa_6_33_0/A dadda_fa_6_33_0/B dadda_fa_6_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_34_0/B dadda_fa_7_33_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_49_0 dadda_fa_3_49_0/A dadda_fa_3_49_0/B dadda_fa_3_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/B dadda_fa_4_49_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2002 U$$84/A1 U$$2048/A2 U$$86/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$2003/A sky130_fd_sc_hd__a22o_1
XU$$2013 U$$2013/A U$$2023/B VGND VGND VPWR VPWR U$$2013/X sky130_fd_sc_hd__xor2_1
XU$$2024 U$$928/A1 U$$2036/A2 _602_/Q U$$2036/B2 VGND VGND VPWR VPWR U$$2025/A sky130_fd_sc_hd__a22o_1
XU$$2035 U$$2035/A U$$2055/A VGND VGND VPWR VPWR U$$2035/X sky130_fd_sc_hd__xor2_1
XU$$2046 U$$950/A1 U$$2052/A2 U$$952/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2047/A sky130_fd_sc_hd__a22o_1
XU$$1301 U$$68/A1 U$$1341/A2 U$$68/B1 U$$1341/B2 VGND VGND VPWR VPWR U$$1302/A sky130_fd_sc_hd__a22o_1
XU$$2057 U$$2186/B VGND VGND VPWR VPWR U$$2057/Y sky130_fd_sc_hd__inv_1
XU$$1312 U$$1312/A U$$1369/A VGND VGND VPWR VPWR U$$1312/X sky130_fd_sc_hd__xor2_1
XFILLER_50_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1323 U$$90/A1 U$$1341/A2 U$$92/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1324/A sky130_fd_sc_hd__a22o_1
XU$$2068 U$$2068/A U$$2118/B VGND VGND VPWR VPWR U$$2068/X sky130_fd_sc_hd__xor2_1
XU$$1334 U$$1334/A U$$1336/B VGND VGND VPWR VPWR U$$1334/X sky130_fd_sc_hd__xor2_1
XU$$2079 _560_/Q U$$2117/A2 _561_/Q U$$2117/B2 VGND VGND VPWR VPWR U$$2080/A sky130_fd_sc_hd__a22o_1
XU$$1345 U$$934/A1 U$$1367/A2 U$$936/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1346/A sky130_fd_sc_hd__a22o_1
XU$$1356 U$$1356/A U$$1369/A VGND VGND VPWR VPWR U$$1356/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_114_1 U$$3826/X U$$3959/X VGND VGND VPWR VPWR dadda_fa_4_115_2/B dadda_ha_3_114_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1367 U$$956/A1 U$$1367/A2 U$$1367/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1368/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1378 U$$8/A1 U$$1474/A2 U$$8/B1 U$$1466/B2 VGND VGND VPWR VPWR U$$1379/A sky130_fd_sc_hd__a22o_1
XU$$1389 U$$1389/A U$$1479/B VGND VGND VPWR VPWR U$$1389/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_106_0 dadda_fa_7_106_0/A dadda_fa_7_106_0/B dadda_fa_7_106_0/CIN VGND
+ VGND VPWR VPWR _531_/D _402_/D sky130_fd_sc_hd__fa_2
XFILLER_157_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_10_clk _431_/CLK VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_51_0 input203/X dadda_fa_2_51_0/B dadda_fa_2_51_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_52_0/B dadda_fa_3_51_2/B sky130_fd_sc_hd__fa_2
Xclkbuf_leaf_77_clk _560_/CLK VGND VGND VPWR VPWR _650_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$30 _454_/Q _326_/Q VGND VGND VPWR VPWR final_adder.U$$525/B1 final_adder.U$$652/A
+ sky130_fd_sc_hd__ha_1
XFILLER_54_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$41 _465_/Q _337_/Q VGND VGND VPWR VPWR final_adder.U$$169/B1 final_adder.U$$663/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$52 _476_/Q _348_/Q VGND VGND VPWR VPWR final_adder.U$$547/B1 final_adder.U$$674/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3270 U$$3270/A U$$3270/B VGND VGND VPWR VPWR U$$3270/X sky130_fd_sc_hd__xor2_1
XU$$3281 _613_/Q U$$3155/X U$$4379/A1 U$$3156/X VGND VGND VPWR VPWR U$$3282/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$63 _487_/Q _359_/Q VGND VGND VPWR VPWR final_adder.U$$191/B1 final_adder.U$$685/A
+ sky130_fd_sc_hd__ha_1
XU$$3292 U$$3290/Y _664_/Q _663_/Q U$$3291/X U$$3288/Y VGND VGND VPWR VPWR U$$3292/X
+ sky130_fd_sc_hd__a32o_4
Xfinal_adder.U$$74 _498_/Q _370_/Q VGND VGND VPWR VPWR final_adder.U$$569/B1 final_adder.U$$696/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$85 _509_/Q _381_/Q VGND VGND VPWR VPWR final_adder.U$$213/B1 final_adder.U$$707/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$96 _520_/Q _392_/Q VGND VGND VPWR VPWR final_adder.U$$591/B1 final_adder.U$$718/A
+ sky130_fd_sc_hd__ha_2
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2580 _605_/Q U$$2470/X _606_/Q U$$2471/X VGND VGND VPWR VPWR U$$2581/A sky130_fd_sc_hd__a22o_1
XU$$2591 U$$2591/A U$$2603/A VGND VGND VPWR VPWR U$$2591/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1890 U$$1890/A U$$1904/B VGND VGND VPWR VPWR U$$1890/X sky130_fd_sc_hd__xor2_1
XFILLER_148_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_80_2 dadda_fa_4_80_2/A dadda_fa_4_80_2/B dadda_fa_4_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/CIN dadda_fa_5_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_73_1 dadda_fa_4_73_1/A dadda_fa_4_73_1/B dadda_fa_4_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/B dadda_fa_5_73_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_89_1 U$$2180/X U$$2313/X U$$2446/X VGND VGND VPWR VPWR dadda_fa_2_90_4/A
+ dadda_fa_2_89_5/B sky130_fd_sc_hd__fa_2
XFILLER_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_50_0 dadda_fa_7_50_0/A dadda_fa_7_50_0/B dadda_fa_7_50_0/CIN VGND VGND
+ VPWR VPWR _475_/D _346_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_66_0 dadda_fa_4_66_0/A dadda_fa_4_66_0/B dadda_fa_4_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/A dadda_fa_5_66_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_68_clk _560_/CLK VGND VGND VPWR VPWR _678_/CLK sky130_fd_sc_hd__clkbuf_16
Xfinal_adder.U$$531 final_adder.U$$658/A final_adder.U$$658/B final_adder.U$$531/B1
+ VGND VGND VPWR VPWR final_adder.U$$659/B sky130_fd_sc_hd__a21o_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_630_ _642_/CLK _630_/D VGND VGND VPWR VPWR _630_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$553 final_adder.U$$680/A final_adder.U$$680/B final_adder.U$$553/B1
+ VGND VGND VPWR VPWR final_adder.U$$681/B sky130_fd_sc_hd__a21o_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$403 U$$403/A _621_/Q VGND VGND VPWR VPWR U$$403/X sky130_fd_sc_hd__xor2_1
XFILLER_85_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$575 final_adder.U$$702/A final_adder.U$$702/B final_adder.U$$575/B1
+ VGND VGND VPWR VPWR final_adder.U$$703/B sky130_fd_sc_hd__a21o_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$414 _623_/Q U$$414/B VGND VGND VPWR VPWR U$$414/X sky130_fd_sc_hd__and2_1
XFILLER_85_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$425 U$$12/B1 U$$545/A2 U$$16/A1 U$$416/X VGND VGND VPWR VPWR U$$426/A sky130_fd_sc_hd__a22o_1
X_561_ _639_/CLK _561_/D VGND VGND VPWR VPWR _561_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$597 final_adder.U$$724/A final_adder.U$$724/B final_adder.U$$597/B1
+ VGND VGND VPWR VPWR final_adder.U$$725/B sky130_fd_sc_hd__a21o_1
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$436 U$$436/A U$$530/B VGND VGND VPWR VPWR U$$436/X sky130_fd_sc_hd__xor2_1
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$447 U$$36/A1 U$$491/A2 U$$38/A1 U$$416/X VGND VGND VPWR VPWR U$$448/A sky130_fd_sc_hd__a22o_1
XU$$458 U$$458/A U$$530/B VGND VGND VPWR VPWR U$$458/X sky130_fd_sc_hd__xor2_1
XU$$469 U$$58/A1 U$$545/A2 U$$60/A1 U$$416/X VGND VGND VPWR VPWR U$$470/A sky130_fd_sc_hd__a22o_1
X_492_ _492_/CLK _492_/D VGND VGND VPWR VPWR _492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_711__763 VGND VGND VPWR VPWR _711__763/HI U$$1093/B1 sky130_fd_sc_hd__conb_1
XFILLER_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_clk _536_/CLK VGND VGND VPWR VPWR _594_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$970 U$$970/A U$$998/B VGND VGND VPWR VPWR U$$970/X sky130_fd_sc_hd__xor2_1
XFILLER_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$981 _559_/Q U$$999/A2 U$$983/A1 U$$999/B2 VGND VGND VPWR VPWR U$$982/A sky130_fd_sc_hd__a22o_1
XU$$1120 U$$983/A1 U$$1200/A2 U$$26/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1121/A sky130_fd_sc_hd__a22o_1
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1131 U$$1131/A U$$1189/B VGND VGND VPWR VPWR U$$1131/X sky130_fd_sc_hd__xor2_1
XU$$992 U$$992/A U$$992/B VGND VGND VPWR VPWR U$$992/X sky130_fd_sc_hd__xor2_1
XFILLER_44_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1142 U$$868/A1 U$$1200/A2 U$$48/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1143/A sky130_fd_sc_hd__a22o_1
XFILLER_188_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1153 U$$1153/A U$$1189/B VGND VGND VPWR VPWR U$$1153/X sky130_fd_sc_hd__xor2_1
XU$$1164 U$$68/A1 U$$1200/A2 U$$68/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1165/A sky130_fd_sc_hd__a22o_1
XFILLER_149_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1175 U$$1175/A U$$1232/A VGND VGND VPWR VPWR U$$1175/X sky130_fd_sc_hd__xor2_1
XFILLER_176_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1186 U$$90/A1 U$$1200/A2 U$$92/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1187/A sky130_fd_sc_hd__a22o_1
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1197 U$$1197/A _633_/Q VGND VGND VPWR VPWR U$$1197/X sky130_fd_sc_hd__xor2_1
XFILLER_54_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_90_1 dadda_fa_5_90_1/A dadda_fa_5_90_1/B dadda_fa_5_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/B dadda_fa_7_90_0/A sky130_fd_sc_hd__fa_1
XFILLER_145_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_83_0 dadda_fa_5_83_0/A dadda_fa_5_83_0/B dadda_fa_5_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/A dadda_fa_6_83_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_99_0 U$$2465/Y U$$2599/X U$$2732/X VGND VGND VPWR VPWR dadda_fa_3_100_1/A
+ dadda_fa_3_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_75_7 U$$4413/X input229/X dadda_fa_1_75_7/CIN VGND VGND VPWR VPWR dadda_fa_2_76_2/CIN
+ dadda_fa_2_75_5/CIN sky130_fd_sc_hd__fa_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_6 dadda_fa_1_68_6/A dadda_fa_1_68_6/B dadda_fa_1_68_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/B dadda_fa_2_68_5/B sky130_fd_sc_hd__fa_2
XFILLER_105_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_701__921 VGND VGND VPWR VPWR _701__921/HI _701__921/LO sky130_fd_sc_hd__conb_1
XFILLER_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_98_0 dadda_fa_7_98_0/A dadda_fa_7_98_0/B dadda_fa_7_98_0/CIN VGND VGND
+ VPWR VPWR _523_/D _394_/D sky130_fd_sc_hd__fa_2
XFILLER_139_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_113_0 dadda_fa_6_113_0/A dadda_fa_6_113_0/B dadda_fa_6_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_114_0/B dadda_fa_7_113_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$361 final_adder.U$$360/A final_adder.U$$337/X final_adder.U$$339/X
+ VGND VGND VPWR VPWR final_adder.U$$361/X sky130_fd_sc_hd__a21o_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$200 U$$200/A U$$274/A VGND VGND VPWR VPWR U$$200/X sky130_fd_sc_hd__xor2_1
XFILLER_73_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_613_ _677_/CLK _613_/D VGND VGND VPWR VPWR _613_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$372 final_adder.U$$372/A final_adder.U$$372/B VGND VGND VPWR VPWR
+ final_adder.U$$372/X sky130_fd_sc_hd__and2_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$211 U$$759/A1 U$$141/X U$$759/B1 U$$142/X VGND VGND VPWR VPWR U$$212/A sky130_fd_sc_hd__a22o_1
XFILLER_40_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$383 final_adder.U$$372/X final_adder.U$$686/B final_adder.U$$373/X
+ VGND VGND VPWR VPWR final_adder.U$$718/B sky130_fd_sc_hd__a21o_2
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$222 U$$222/A U$$274/A VGND VGND VPWR VPWR U$$222/X sky130_fd_sc_hd__xor2_1
XFILLER_73_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_33_3 dadda_fa_3_33_3/A dadda_fa_3_33_3/B dadda_fa_3_33_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/B dadda_fa_4_33_2/CIN sky130_fd_sc_hd__fa_2
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$233 U$$94/B1 U$$141/X U$$98/A1 U$$142/X VGND VGND VPWR VPWR U$$234/A sky130_fd_sc_hd__a22o_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$244 U$$244/A U$$262/B VGND VGND VPWR VPWR U$$244/X sky130_fd_sc_hd__xor2_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$255 U$$940/A1 U$$141/X U$$942/A1 U$$142/X VGND VGND VPWR VPWR U$$256/A sky130_fd_sc_hd__a22o_1
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_544_ _678_/CLK _544_/D VGND VGND VPWR VPWR _544_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_2 U$$1918/A input175/X dadda_fa_3_26_2/CIN VGND VGND VPWR VPWR dadda_fa_4_27_1/A
+ dadda_fa_4_26_2/B sky130_fd_sc_hd__fa_2
XU$$266 U$$266/A _619_/Q VGND VGND VPWR VPWR U$$266/X sky130_fd_sc_hd__xor2_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$277 _621_/Q U$$277/B VGND VGND VPWR VPWR U$$277/X sky130_fd_sc_hd__and2_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$288 U$$12/B1 U$$278/X U$$16/A1 U$$279/X VGND VGND VPWR VPWR U$$289/A sky130_fd_sc_hd__a22o_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_19_1 U$$444/X U$$577/X U$$710/X VGND VGND VPWR VPWR dadda_fa_4_20_1/A
+ dadda_fa_4_19_2/B sky130_fd_sc_hd__fa_2
XU$$299 U$$299/A U$$357/B VGND VGND VPWR VPWR U$$299/X sky130_fd_sc_hd__xor2_1
XFILLER_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_475_ _483_/CLK _475_/D VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$5 U$$3/B U$$5/A2 U$$1/A U$$0/Y VGND VGND VPWR VPWR U$$5/X sky130_fd_sc_hd__a22o_4
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput308 _198_/Q VGND VGND VPWR VPWR o[30] sky130_fd_sc_hd__buf_2
XFILLER_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput319 _208_/Q VGND VGND VPWR VPWR o[40] sky130_fd_sc_hd__buf_2
XFILLER_142_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_78_5 dadda_fa_2_78_5/A dadda_fa_2_78_5/B dadda_fa_2_78_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_2/A dadda_fa_4_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_108_1 dadda_fa_5_108_1/A dadda_fa_5_108_1/B dadda_fa_5_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/B dadda_fa_7_108_0/A sky130_fd_sc_hd__fa_2
XFILLER_191_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_5 U$$3093/X U$$3226/X U$$3359/X VGND VGND VPWR VPWR dadda_fa_2_81_2/B
+ dadda_fa_2_80_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_73_4 U$$3478/X U$$3611/X U$$3744/X VGND VGND VPWR VPWR dadda_fa_2_74_1/CIN
+ dadda_fa_2_73_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_66_3 U$$3730/X U$$3863/X U$$3996/X VGND VGND VPWR VPWR dadda_fa_2_67_1/B
+ dadda_fa_2_66_4/B sky130_fd_sc_hd__fa_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_43_2 dadda_fa_4_43_2/A dadda_fa_4_43_2/B dadda_fa_4_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/CIN dadda_fa_5_43_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_59_2 U$$2386/X U$$2519/X U$$2652/X VGND VGND VPWR VPWR dadda_fa_2_60_1/A
+ dadda_fa_2_59_4/A sky130_fd_sc_hd__fa_1
XFILLER_6_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_36_1 dadda_fa_4_36_1/A dadda_fa_4_36_1/B dadda_fa_4_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/B dadda_fa_5_36_1/B sky130_fd_sc_hd__fa_1
XFILLER_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_13_0 dadda_fa_7_13_0/A dadda_fa_7_13_0/B dadda_fa_7_13_0/CIN VGND VGND
+ VPWR VPWR _438_/D _309_/D sky130_fd_sc_hd__fa_2
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_0 dadda_fa_4_29_0/A dadda_fa_4_29_0/B dadda_fa_4_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/A dadda_fa_5_29_1/A sky130_fd_sc_hd__fa_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_260_ _379_/CLK _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_191_ _333_/CLK _191_/D VGND VGND VPWR VPWR _191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4504 U$$4504/A1 U$$4388/X U$$4506/A1 U$$4389/X VGND VGND VPWR VPWR U$$4505/A sky130_fd_sc_hd__a22o_1
XU$$4515 U$$4515/A U$$4515/B VGND VGND VPWR VPWR U$$4515/X sky130_fd_sc_hd__xor2_2
X_782__834 VGND VGND VPWR VPWR _782__834/HI U$$4409/B sky130_fd_sc_hd__conb_1
Xdadda_fa_0_61_2 U$$927/X U$$1060/X U$$1193/X VGND VGND VPWR VPWR dadda_fa_1_62_6/B
+ dadda_fa_1_61_8/B sky130_fd_sc_hd__fa_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3803 U$$787/B1 U$$3703/X U$$654/A1 U$$3704/X VGND VGND VPWR VPWR U$$3804/A sky130_fd_sc_hd__a22o_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3814 U$$3814/A U$$3835/A VGND VGND VPWR VPWR U$$3814/X sky130_fd_sc_hd__xor2_1
XU$$18 U$$18/A1 U$$4/X U$$20/A1 U$$5/X VGND VGND VPWR VPWR U$$19/A sky130_fd_sc_hd__a22o_1
XFILLER_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$29 U$$29/A U$$89/B VGND VGND VPWR VPWR U$$29/X sky130_fd_sc_hd__xor2_1
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3825 _611_/Q U$$3703/X U$$539/A1 U$$3704/X VGND VGND VPWR VPWR U$$3826/A sky130_fd_sc_hd__a22o_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3836 _671_/Q VGND VGND VPWR VPWR U$$3836/Y sky130_fd_sc_hd__inv_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_0 U$$1931/X U$$2064/X input181/X VGND VGND VPWR VPWR dadda_fa_4_32_0/B
+ dadda_fa_4_31_1/CIN sky130_fd_sc_hd__fa_2
XU$$3847 U$$3847/A U$$3893/B VGND VGND VPWR VPWR U$$3847/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$180 final_adder.U$$675/A final_adder.U$$674/A VGND VGND VPWR VPWR
+ final_adder.U$$282/B sky130_fd_sc_hd__and2_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3858 _559_/Q U$$3912/A2 _560_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3859/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$191 final_adder.U$$685/A final_adder.U$$557/B1 final_adder.U$$191/B1
+ VGND VGND VPWR VPWR final_adder.U$$191/X sky130_fd_sc_hd__a21o_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3869 U$$3869/A U$$3929/B VGND VGND VPWR VPWR U$$3869/X sky130_fd_sc_hd__xor2_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_823__875 VGND VGND VPWR VPWR _823__875/HI U$$4491/B sky130_fd_sc_hd__conb_1
XFILLER_72_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_527_ _527_/CLK _527_/D VGND VGND VPWR VPWR _527_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_458_ _458_/CLK _458_/D VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_389_ _535_/CLK _389_/D VGND VGND VPWR VPWR _389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_90_4 dadda_fa_2_90_4/A dadda_fa_2_90_4/B dadda_fa_2_90_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_1/CIN dadda_fa_3_90_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_83_3 dadda_fa_2_83_3/A dadda_fa_2_83_3/B dadda_fa_2_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/B dadda_fa_3_83_3/B sky130_fd_sc_hd__fa_1
XFILLER_141_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_76_2 dadda_fa_2_76_2/A dadda_fa_2_76_2/B dadda_fa_2_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/A dadda_fa_3_76_3/A sky130_fd_sc_hd__fa_2
Xdadda_fa_5_53_1 dadda_fa_5_53_1/A dadda_fa_5_53_1/B dadda_fa_5_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/B dadda_fa_7_53_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_69_1 dadda_fa_2_69_1/A dadda_fa_2_69_1/B dadda_fa_2_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/CIN dadda_fa_3_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_46_0 dadda_fa_5_46_0/A dadda_fa_5_46_0/B dadda_fa_5_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/A dadda_fa_6_46_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_120_0 U$$4503/X input152/X dadda_fa_5_120_0/CIN VGND VGND VPWR VPWR dadda_fa_6_121_0/A
+ dadda_fa_6_120_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_71_1 U$$2543/X U$$2676/X U$$2809/X VGND VGND VPWR VPWR dadda_fa_2_72_0/CIN
+ dadda_fa_2_71_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_160_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_766__818 VGND VGND VPWR VPWR _766__818/HI U$$4381/B1 sky130_fd_sc_hd__conb_1
XFILLER_8_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_64_0 U$$2529/X U$$2662/X U$$2795/X VGND VGND VPWR VPWR dadda_fa_2_65_0/B
+ dadda_fa_2_64_3/B sky130_fd_sc_hd__fa_1
XFILLER_143_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_807__859 VGND VGND VPWR VPWR _807__859/HI U$$4459/B sky130_fd_sc_hd__conb_1
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2409 _588_/Q U$$2421/A2 _589_/Q U$$2421/B2 VGND VGND VPWR VPWR U$$2410/A sky130_fd_sc_hd__a22o_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1708 U$$3900/A1 U$$1726/A2 U$$3489/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1709/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1719 U$$1719/A U$$1739/B VGND VGND VPWR VPWR U$$1719/X sky130_fd_sc_hd__xor2_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _452_/CLK _312_/D VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_243_ _501_/CLK _243_/D VGND VGND VPWR VPWR _243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 a[25] VGND VGND VPWR VPWR _641_/D sky130_fd_sc_hd__clkbuf_2
X_174_ _462_/CLK _174_/D VGND VGND VPWR VPWR _174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 a[35] VGND VGND VPWR VPWR _651_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_182_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_93_2 dadda_fa_3_93_2/A dadda_fa_3_93_2/B dadda_fa_3_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/A dadda_fa_4_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_183_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_86_1 dadda_fa_3_86_1/A dadda_fa_3_86_1/B dadda_fa_3_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/CIN dadda_fa_4_86_2/A sky130_fd_sc_hd__fa_2
XFILLER_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_63_0 dadda_fa_6_63_0/A dadda_fa_6_63_0/B dadda_fa_6_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_64_0/B dadda_fa_7_63_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_97_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_79_0 dadda_fa_3_79_0/A dadda_fa_3_79_0/B dadda_fa_3_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/B dadda_fa_4_79_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_53_0 U$$113/X U$$246/X VGND VGND VPWR VPWR dadda_fa_1_54_8/B dadda_fa_2_53_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater608 _619_/Q VGND VGND VPWR VPWR U$$262/B sky130_fd_sc_hd__buf_12
XFILLER_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4301 _575_/Q U$$4251/X U$$4303/A1 U$$4252/X VGND VGND VPWR VPWR U$$4302/A sky130_fd_sc_hd__a22o_1
Xrepeater619 _612_/Q VGND VGND VPWR VPWR U$$950/A1 sky130_fd_sc_hd__buf_12
XU$$4312 U$$4312/A U$$4384/A VGND VGND VPWR VPWR U$$4312/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4323 U$$759/B1 U$$4377/A2 U$$78/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4324/A sky130_fd_sc_hd__a22o_1
XU$$4334 U$$4334/A _679_/Q VGND VGND VPWR VPWR U$$4334/X sky130_fd_sc_hd__xor2_1
XU$$4345 U$$98/A1 U$$4381/A2 U$$4484/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4346/A sky130_fd_sc_hd__a22o_1
XU$$3600 U$$4285/A1 U$$3624/A2 U$$4424/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3601/A
+ sky130_fd_sc_hd__a22o_1
XU$$3611 U$$3611/A U$$3699/A VGND VGND VPWR VPWR U$$3611/X sky130_fd_sc_hd__xor2_1
XU$$4356 U$$4356/A _679_/Q VGND VGND VPWR VPWR U$$4356/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_1 U$$4360/X U$$4493/X input146/X VGND VGND VPWR VPWR dadda_fa_5_116_0/B
+ dadda_fa_5_115_1/B sky130_fd_sc_hd__fa_1
XU$$4367 U$$4504/A1 U$$4377/A2 U$$4506/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4368/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3622 U$$4170/A1 U$$3624/A2 U$$3624/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3623/A
+ sky130_fd_sc_hd__a22o_1
XU$$3633 U$$3633/A U$$3699/A VGND VGND VPWR VPWR U$$3633/X sky130_fd_sc_hd__xor2_1
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4378 U$$4378/A U$$4384/A VGND VGND VPWR VPWR U$$4378/X sky130_fd_sc_hd__xor2_1
XU$$3644 _589_/Q U$$3668/A2 _590_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3645/A sky130_fd_sc_hd__a22o_1
XU$$4389 U$$4387/B U$$4384/A U$$4389/B1 U$$4384/Y VGND VGND VPWR VPWR U$$4389/X sky130_fd_sc_hd__a22o_4
XFILLER_34_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2910 U$$2910/A U$$2996/B VGND VGND VPWR VPWR U$$2910/X sky130_fd_sc_hd__xor2_1
XU$$3655 U$$3655/A U$$3699/A VGND VGND VPWR VPWR U$$3655/X sky130_fd_sc_hd__xor2_1
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_108_0 dadda_fa_4_108_0/A dadda_fa_4_108_0/B dadda_fa_4_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/A dadda_fa_5_108_1/A sky130_fd_sc_hd__fa_1
XU$$3666 _600_/Q U$$3668/A2 _601_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3667/A sky130_fd_sc_hd__a22o_1
XU$$2921 U$$4289/B1 U$$2975/A2 U$$4291/B1 U$$2975/B2 VGND VGND VPWR VPWR U$$2922/A
+ sky130_fd_sc_hd__a22o_1
XU$$3677 U$$3677/A U$$3698/A VGND VGND VPWR VPWR U$$3677/X sky130_fd_sc_hd__xor2_1
XU$$2932 U$$2932/A U$$2996/B VGND VGND VPWR VPWR U$$2932/X sky130_fd_sc_hd__xor2_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2943 _581_/Q U$$2881/X U$$4178/A1 U$$2882/X VGND VGND VPWR VPWR U$$2944/A sky130_fd_sc_hd__a22o_1
XU$$3688 U$$4510/A1 U$$3566/X U$$539/A1 U$$3567/X VGND VGND VPWR VPWR U$$3689/A sky130_fd_sc_hd__a22o_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2954 U$$2954/A U$$2960/B VGND VGND VPWR VPWR U$$2954/X sky130_fd_sc_hd__xor2_1
XFILLER_18_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3699 U$$3699/A VGND VGND VPWR VPWR U$$3699/Y sky130_fd_sc_hd__inv_1
XU$$2965 U$$4335/A1 U$$2881/X _593_/Q U$$2882/X VGND VGND VPWR VPWR U$$2966/A sky130_fd_sc_hd__a22o_1
XU$$2976 U$$2976/A _659_/Q VGND VGND VPWR VPWR U$$2976/X sky130_fd_sc_hd__xor2_1
XU$$2987 U$$932/A1 U$$3009/A2 U$$934/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2988/A sky130_fd_sc_hd__a22o_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2998 U$$2998/A U$$3004/B VGND VGND VPWR VPWR U$$2998/X sky130_fd_sc_hd__xor2_1
XFILLER_33_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_81_0 U$$4425/X input236/X dadda_fa_2_81_0/CIN VGND VGND VPWR VPWR dadda_fa_3_82_0/B
+ dadda_fa_3_81_2/B sky130_fd_sc_hd__fa_2
XFILLER_138_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_51_8 U$$3301/X U$$3434/X VGND VGND VPWR VPWR dadda_fa_2_52_3/A dadda_fa_3_51_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_130_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_50_6 U$$2501/X U$$2634/X U$$2767/X VGND VGND VPWR VPWR dadda_fa_2_51_2/B
+ dadda_fa_2_50_5/B sky130_fd_sc_hd__fa_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_2_0 U$$242/B input179/X dadda_ha_6_2_0/SUM VGND VGND VPWR VPWR _427_/D
+ _298_/D sky130_fd_sc_hd__fa_1
XFILLER_97_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_80_0 dadda_fa_7_80_0/A dadda_fa_7_80_0/B dadda_fa_7_80_0/CIN VGND VGND
+ VPWR VPWR _505_/D _376_/D sky130_fd_sc_hd__fa_1
XFILLER_192_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_96_0 dadda_fa_4_96_0/A dadda_fa_4_96_0/B dadda_fa_4_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/A dadda_fa_5_96_1/A sky130_fd_sc_hd__fa_2
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2206 U$$14/A1 U$$2270/A2 U$$14/B1 U$$2286/B2 VGND VGND VPWR VPWR U$$2207/A sky130_fd_sc_hd__a22o_1
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2217 U$$2217/A U$$2257/B VGND VGND VPWR VPWR U$$2217/X sky130_fd_sc_hd__xor2_1
XU$$2228 U$$36/A1 U$$2196/X _567_/Q U$$2197/X VGND VGND VPWR VPWR U$$2229/A sky130_fd_sc_hd__a22o_1
XU$$2239 U$$2239/A U$$2257/B VGND VGND VPWR VPWR U$$2239/X sky130_fd_sc_hd__xor2_1
XU$$1505 U$$1505/A U$$1505/B VGND VGND VPWR VPWR U$$1505/X sky130_fd_sc_hd__xor2_1
XU$$1516 U$$1516/A U$$1614/B VGND VGND VPWR VPWR U$$1516/X sky130_fd_sc_hd__xor2_1
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1527 U$$842/A1 U$$1511/X U$$22/A1 U$$1512/X VGND VGND VPWR VPWR U$$1528/A sky130_fd_sc_hd__a22o_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1538 U$$1538/A U$$1580/B VGND VGND VPWR VPWR U$$1538/X sky130_fd_sc_hd__xor2_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1549 U$$3876/B1 U$$1591/A2 U$$4291/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1550/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ _474_/CLK _226_/D VGND VGND VPWR VPWR _226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_788__840 VGND VGND VPWR VPWR _788__840/HI U$$4421/B sky130_fd_sc_hd__conb_1
XFILLER_3_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_60_5 dadda_fa_2_60_5/A dadda_fa_2_60_5/B dadda_fa_2_60_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_2/A dadda_fa_4_60_0/A sky130_fd_sc_hd__fa_2
XFILLER_66_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater405 U$$3678/A2 VGND VGND VPWR VPWR U$$3624/A2 sky130_fd_sc_hd__buf_12
Xrepeater416 U$$2881/X VGND VGND VPWR VPWR U$$2975/A2 sky130_fd_sc_hd__buf_12
Xrepeater427 U$$2333/X VGND VGND VPWR VPWR U$$2463/A2 sky130_fd_sc_hd__buf_12
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_829__881 VGND VGND VPWR VPWR _829__881/HI U$$4503/B sky130_fd_sc_hd__conb_1
XFILLER_66_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_53_4 dadda_fa_2_53_4/A dadda_fa_2_53_4/B dadda_fa_2_53_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/CIN dadda_fa_3_53_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater438 U$$1785/X VGND VGND VPWR VPWR U$$1897/A2 sky130_fd_sc_hd__buf_12
XU$$4120 _553_/Q U$$4114/X U$$4122/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4121/A sky130_fd_sc_hd__a22o_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater449 U$$1237/X VGND VGND VPWR VPWR U$$1367/A2 sky130_fd_sc_hd__buf_12
XU$$4131 U$$4131/A _677_/Q VGND VGND VPWR VPWR U$$4131/X sky130_fd_sc_hd__xor2_1
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4142 _564_/Q U$$4198/A2 _565_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4143/A sky130_fd_sc_hd__a22o_1
XU$$4153 U$$4153/A U$$4197/B VGND VGND VPWR VPWR U$$4153/X sky130_fd_sc_hd__xor2_1
XFILLER_65_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_46_3 dadda_fa_2_46_3/A dadda_fa_2_46_3/B dadda_fa_2_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/B dadda_fa_3_46_3/B sky130_fd_sc_hd__fa_2
XU$$4164 U$$4438/A1 U$$4198/A2 U$$56/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4165/A sky130_fd_sc_hd__a22o_1
XU$$3430 U$$3428/B _665_/Q _666_/Q U$$3425/Y VGND VGND VPWR VPWR U$$3430/X sky130_fd_sc_hd__a22o_4
XU$$4175 U$$4175/A U$$4247/A VGND VGND VPWR VPWR U$$4175/X sky130_fd_sc_hd__xor2_1
XU$$3441 U$$16/A1 U$$3429/X U$$975/B1 U$$3430/X VGND VGND VPWR VPWR U$$3442/A sky130_fd_sc_hd__a22o_1
XU$$4186 _586_/Q U$$4114/X _587_/Q U$$4115/X VGND VGND VPWR VPWR U$$4187/A sky130_fd_sc_hd__a22o_1
XU$$4197 U$$4197/A U$$4197/B VGND VGND VPWR VPWR U$$4197/X sky130_fd_sc_hd__xor2_1
XU$$3452 U$$3452/A U$$3496/B VGND VGND VPWR VPWR U$$3452/X sky130_fd_sc_hd__xor2_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_39_2 U$$1947/X U$$2080/X U$$2213/X VGND VGND VPWR VPWR dadda_fa_3_40_1/A
+ dadda_fa_3_39_3/A sky130_fd_sc_hd__fa_1
XU$$3463 _567_/Q U$$3545/A2 U$$4424/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3464/A sky130_fd_sc_hd__a22o_1
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3474 U$$3474/A U$$3496/B VGND VGND VPWR VPWR U$$3474/X sky130_fd_sc_hd__xor2_1
XU$$3485 U$$4170/A1 U$$3545/A2 U$$3624/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3486/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_16_1 dadda_fa_5_16_1/A dadda_fa_5_16_1/B dadda_fa_5_16_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/B dadda_fa_7_16_0/A sky130_fd_sc_hd__fa_2
XU$$2740 _655_/Q VGND VGND VPWR VPWR U$$2740/Y sky130_fd_sc_hd__inv_1
XU$$2751 U$$2751/A U$$2797/B VGND VGND VPWR VPWR U$$2751/X sky130_fd_sc_hd__xor2_1
XU$$3496 U$$3496/A U$$3496/B VGND VGND VPWR VPWR U$$3496/X sky130_fd_sc_hd__xor2_1
XU$$2762 U$$979/B1 U$$2796/A2 U$$983/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2763/A sky130_fd_sc_hd__a22o_1
XU$$2773 U$$2773/A U$$2839/B VGND VGND VPWR VPWR U$$2773/X sky130_fd_sc_hd__xor2_1
XFILLER_179_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2784 U$$4289/B1 U$$2870/A2 U$$4291/B1 U$$2834/B2 VGND VGND VPWR VPWR U$$2785/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2795 U$$2795/A U$$2797/B VGND VGND VPWR VPWR U$$2795/X sky130_fd_sc_hd__xor2_1
XFILLER_22_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_42_4 U$$1687/X U$$1820/X VGND VGND VPWR VPWR dadda_fa_2_43_4/B dadda_fa_3_42_0/A
+ sky130_fd_sc_hd__ha_2
Xinput208 c[56] VGND VGND VPWR VPWR input208/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput219 c[66] VGND VGND VPWR VPWR input219/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfinal_adder.U$$702 final_adder.U$$702/A final_adder.U$$702/B VGND VGND VPWR VPWR
+ _248_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$713 final_adder.U$$713/A final_adder.U$$713/B VGND VGND VPWR VPWR
+ _259_/D sky130_fd_sc_hd__xor2_2
XFILLER_151_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$724 final_adder.U$$724/A final_adder.U$$724/B VGND VGND VPWR VPWR
+ _270_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_4_12_2 U$$829/X U$$903/B VGND VGND VPWR VPWR dadda_fa_5_13_0/CIN dadda_ha_4_12_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_84_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$735 final_adder.U$$735/A final_adder.U$$735/B VGND VGND VPWR VPWR
+ _281_/D sky130_fd_sc_hd__xor2_1
XFILLER_112_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$746 final_adder.U$$746/A final_adder.U$$746/B VGND VGND VPWR VPWR
+ _292_/D sky130_fd_sc_hd__xor2_1
XFILLER_151_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$607 U$$607/A U$$661/B VGND VGND VPWR VPWR U$$607/X sky130_fd_sc_hd__xor2_1
XFILLER_72_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$618 U$$70/A1 U$$626/A2 U$$70/B1 U$$553/X VGND VGND VPWR VPWR U$$619/A sky130_fd_sc_hd__a22o_1
XFILLER_99_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_41_2 U$$887/X U$$1020/X U$$1153/X VGND VGND VPWR VPWR dadda_fa_2_42_4/A
+ dadda_fa_2_41_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$629 U$$629/A U$$661/B VGND VGND VPWR VPWR U$$629/X sky130_fd_sc_hd__xor2_1
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_11_0 U$$29/X U$$162/X U$$295/X VGND VGND VPWR VPWR dadda_fa_5_12_0/B dadda_fa_5_11_1/B
+ sky130_fd_sc_hd__fa_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_115_0 U$$3561/Y U$$3695/X U$$3828/X VGND VGND VPWR VPWR dadda_fa_4_116_2/B
+ dadda_fa_4_115_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_192_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_63_3 dadda_fa_3_63_3/A dadda_fa_3_63_3/B dadda_fa_3_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/B dadda_fa_4_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_56_2 dadda_fa_3_56_2/A dadda_fa_3_56_2/B dadda_fa_3_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/A dadda_fa_4_56_2/B sky130_fd_sc_hd__fa_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_49_1 dadda_fa_3_49_1/A dadda_fa_3_49_1/B dadda_fa_3_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/CIN dadda_fa_4_49_2/A sky130_fd_sc_hd__fa_1
XFILLER_63_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_26_0 dadda_fa_6_26_0/A dadda_fa_6_26_0/B dadda_fa_6_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_27_0/B dadda_fa_7_26_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2003 U$$2003/A U$$2023/B VGND VGND VPWR VPWR U$$2003/X sky130_fd_sc_hd__xor2_1
XU$$2014 _596_/Q U$$2036/A2 _597_/Q U$$2036/B2 VGND VGND VPWR VPWR U$$2015/A sky130_fd_sc_hd__a22o_1
XU$$2025 U$$2025/A U$$2055/A VGND VGND VPWR VPWR U$$2025/X sky130_fd_sc_hd__xor2_2
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2036 _607_/Q U$$2036/A2 _608_/Q U$$2036/B2 VGND VGND VPWR VPWR U$$2037/A sky130_fd_sc_hd__a22o_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2047 U$$2047/A _645_/Q VGND VGND VPWR VPWR U$$2047/X sky130_fd_sc_hd__xor2_1
XU$$1302 U$$1302/A U$$1342/B VGND VGND VPWR VPWR U$$1302/X sky130_fd_sc_hd__xor2_1
XU$$1313 U$$902/A1 U$$1367/A2 U$$902/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1314/A sky130_fd_sc_hd__a22o_1
XFILLER_188_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2058 U$$2186/B U$$2058/B VGND VGND VPWR VPWR U$$2058/X sky130_fd_sc_hd__and2_1
XU$$2069 U$$14/A1 U$$2117/A2 U$$14/B1 U$$2117/B2 VGND VGND VPWR VPWR U$$2070/A sky130_fd_sc_hd__a22o_1
XU$$1324 U$$1324/A U$$1342/B VGND VGND VPWR VPWR U$$1324/X sky130_fd_sc_hd__xor2_1
XU$$1335 U$$924/A1 U$$1341/A2 U$$787/B1 U$$1341/B2 VGND VGND VPWR VPWR U$$1336/A sky130_fd_sc_hd__a22o_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1346 U$$1346/A _635_/Q VGND VGND VPWR VPWR U$$1346/X sky130_fd_sc_hd__xor2_1
XFILLER_71_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1357 _610_/Q U$$1367/A2 _611_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1358/A sky130_fd_sc_hd__a22o_1
XFILLER_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1368 U$$1368/A U$$1369/A VGND VGND VPWR VPWR U$$1368/X sky130_fd_sc_hd__xor2_1
XFILLER_71_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1379 U$$1379/A U$$1461/B VGND VGND VPWR VPWR U$$1379/X sky130_fd_sc_hd__xor2_1
XFILLER_176_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ _456_/CLK hold5/X VGND VGND VPWR VPWR _209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_51_1 dadda_fa_2_51_1/A dadda_fa_2_51_1/B dadda_fa_2_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_0/CIN dadda_fa_3_51_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_44_0 U$$2356/X U$$2489/X U$$2622/X VGND VGND VPWR VPWR dadda_fa_3_45_0/B
+ dadda_fa_3_44_2/B sky130_fd_sc_hd__fa_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$20 _444_/Q _316_/Q VGND VGND VPWR VPWR final_adder.U$$515/B1 final_adder.U$$642/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$31 _455_/Q _327_/Q VGND VGND VPWR VPWR final_adder.U$$159/B1 final_adder.U$$653/A
+ sky130_fd_sc_hd__ha_1
XFILLER_81_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3260 U$$3260/A U$$3270/B VGND VGND VPWR VPWR U$$3260/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$42 _466_/Q _338_/Q VGND VGND VPWR VPWR final_adder.U$$537/B1 final_adder.U$$664/A
+ sky130_fd_sc_hd__ha_1
XU$$3271 U$$4504/A1 U$$3155/X U$$4506/A1 U$$3156/X VGND VGND VPWR VPWR U$$3272/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$53 _477_/Q _349_/Q VGND VGND VPWR VPWR final_adder.U$$181/B1 final_adder.U$$675/A
+ sky130_fd_sc_hd__ha_1
XU$$3282 U$$3282/A _663_/Q VGND VGND VPWR VPWR U$$3282/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$64 _488_/Q _360_/Q VGND VGND VPWR VPWR final_adder.U$$559/B1 final_adder.U$$686/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$75 _499_/Q _371_/Q VGND VGND VPWR VPWR final_adder.U$$203/B1 final_adder.U$$697/A
+ sky130_fd_sc_hd__ha_1
XU$$3293 U$$3291/B _663_/Q _664_/Q U$$3288/Y VGND VGND VPWR VPWR U$$3293/X sky130_fd_sc_hd__a22o_4
XFILLER_81_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$86 _510_/Q _382_/Q VGND VGND VPWR VPWR final_adder.U$$581/B1 final_adder.U$$708/A
+ sky130_fd_sc_hd__ha_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2570 U$$787/B1 U$$2470/X _601_/Q U$$2471/X VGND VGND VPWR VPWR U$$2571/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$97 _521_/Q _393_/Q VGND VGND VPWR VPWR final_adder.U$$225/B1 final_adder.U$$719/A
+ sky130_fd_sc_hd__ha_2
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2581 U$$2581/A U$$2603/A VGND VGND VPWR VPWR U$$2581/X sky130_fd_sc_hd__xor2_1
XU$$2592 _611_/Q U$$2470/X _612_/Q U$$2471/X VGND VGND VPWR VPWR U$$2593/A sky130_fd_sc_hd__a22o_1
XFILLER_55_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1880 U$$1880/A U$$1904/B VGND VGND VPWR VPWR U$$1880/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1891 _603_/Q U$$1897/A2 U$$4496/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1892/A sky130_fd_sc_hd__a22o_1
XFILLER_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_73_2 dadda_fa_4_73_2/A dadda_fa_4_73_2/B dadda_fa_4_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/CIN dadda_fa_5_73_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_89_2 U$$2579/X U$$2712/X U$$2845/X VGND VGND VPWR VPWR dadda_fa_2_90_4/B
+ dadda_fa_2_89_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_66_1 dadda_fa_4_66_1/A dadda_fa_4_66_1/B dadda_fa_4_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/B dadda_fa_5_66_1/B sky130_fd_sc_hd__fa_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_43_0 dadda_fa_7_43_0/A dadda_fa_7_43_0/B dadda_fa_7_43_0/CIN VGND VGND
+ VPWR VPWR _468_/D _339_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_59_0 dadda_fa_4_59_0/A dadda_fa_4_59_0/B dadda_fa_4_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/A dadda_fa_5_59_1/A sky130_fd_sc_hd__fa_1
XFILLER_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$521 final_adder.U$$648/A final_adder.U$$648/B final_adder.U$$521/B1
+ VGND VGND VPWR VPWR final_adder.U$$649/B sky130_fd_sc_hd__a21o_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$543 final_adder.U$$670/A final_adder.U$$670/B final_adder.U$$543/B1
+ VGND VGND VPWR VPWR final_adder.U$$671/B sky130_fd_sc_hd__a21o_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$565 final_adder.U$$692/A final_adder.U$$692/B final_adder.U$$565/B1
+ VGND VGND VPWR VPWR final_adder.U$$693/B sky130_fd_sc_hd__a21o_1
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$404 U$$952/A1 U$$278/X U$$952/B1 U$$279/X VGND VGND VPWR VPWR U$$405/A sky130_fd_sc_hd__a22o_1
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$415 U$$413/Y _622_/Q _621_/Q U$$414/X U$$411/Y VGND VGND VPWR VPWR U$$415/X sky130_fd_sc_hd__a32o_4
X_560_ _560_/CLK _560_/D VGND VGND VPWR VPWR _560_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$587 final_adder.U$$714/A final_adder.U$$714/B final_adder.U$$587/B1
+ VGND VGND VPWR VPWR final_adder.U$$715/B sky130_fd_sc_hd__a21o_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$426 U$$426/A _623_/Q VGND VGND VPWR VPWR U$$426/X sky130_fd_sc_hd__xor2_1
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$437 U$$26/A1 U$$491/A2 U$$987/A1 U$$416/X VGND VGND VPWR VPWR U$$438/A sky130_fd_sc_hd__a22o_1
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$448 U$$448/A U$$547/A VGND VGND VPWR VPWR U$$448/X sky130_fd_sc_hd__xor2_1
XU$$459 _572_/Q U$$491/A2 U$$735/A1 U$$416/X VGND VGND VPWR VPWR U$$460/A sky130_fd_sc_hd__a22o_1
X_491_ _492_/CLK _491_/D VGND VGND VPWR VPWR _491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_61_0 dadda_fa_3_61_0/A dadda_fa_3_61_0/B dadda_fa_3_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/B dadda_fa_4_61_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_77_0 U$$958/Y U$$1092/X U$$1225/X VGND VGND VPWR VPWR dadda_fa_1_78_8/CIN
+ dadda_fa_2_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$960 _630_/Q VGND VGND VPWR VPWR U$$962/B sky130_fd_sc_hd__inv_1
Xdadda_ha_4_8_0 U$$23/X U$$156/X VGND VGND VPWR VPWR dadda_fa_5_9_1/B dadda_ha_4_8_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$971 U$$971/A1 U$$963/X U$$12/B1 U$$999/B2 VGND VGND VPWR VPWR U$$972/A sky130_fd_sc_hd__a22o_1
XU$$1110 U$$12/B1 U$$1200/A2 U$$14/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1111/A sky130_fd_sc_hd__a22o_1
XFILLER_90_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$982 U$$982/A U$$992/B VGND VGND VPWR VPWR U$$982/X sky130_fd_sc_hd__xor2_1
XU$$1121 U$$1121/A U$$1189/B VGND VGND VPWR VPWR U$$1121/X sky130_fd_sc_hd__xor2_1
XU$$1132 U$$36/A1 U$$1200/A2 U$$38/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1133/A sky130_fd_sc_hd__a22o_1
XU$$993 U$$34/A1 U$$963/X U$$36/A1 U$$999/B2 VGND VGND VPWR VPWR U$$994/A sky130_fd_sc_hd__a22o_1
XU$$1143 U$$1143/A U$$1167/B VGND VGND VPWR VPWR U$$1143/X sky130_fd_sc_hd__xor2_1
XU$$1154 U$$58/A1 U$$1200/A2 U$$60/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1155/A sky130_fd_sc_hd__a22o_1
XU$$1165 U$$1165/A U$$1167/B VGND VGND VPWR VPWR U$$1165/X sky130_fd_sc_hd__xor2_1
XU$$1176 U$$902/A1 U$$1218/A2 U$$902/B1 U$$1218/B2 VGND VGND VPWR VPWR U$$1177/A sky130_fd_sc_hd__a22o_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1187 U$$1187/A U$$1189/B VGND VGND VPWR VPWR U$$1187/X sky130_fd_sc_hd__xor2_1
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1198 U$$924/A1 U$$1200/A2 U$$787/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1199/A sky130_fd_sc_hd__a22o_1
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_83_1 dadda_fa_5_83_1/A dadda_fa_5_83_1/B dadda_fa_5_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/B dadda_fa_7_83_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_99_1 U$$2865/X U$$2998/X U$$3131/X VGND VGND VPWR VPWR dadda_fa_3_100_1/B
+ dadda_fa_3_99_3/A sky130_fd_sc_hd__fa_1
XFILLER_116_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_76_0 dadda_fa_5_76_0/A dadda_fa_5_76_0/B dadda_fa_5_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/A dadda_fa_6_76_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_75_8 dadda_fa_1_75_8/A dadda_fa_1_75_8/B dadda_fa_1_75_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_76_3/A dadda_fa_3_75_0/A sky130_fd_sc_hd__fa_2
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_7 dadda_fa_1_68_7/A dadda_fa_1_68_7/B dadda_fa_1_68_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/CIN dadda_fa_2_68_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3090 U$$76/A1 U$$3090/A2 U$$78/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3091/A sky130_fd_sc_hd__a22o_1
XFILLER_35_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_734__786 VGND VGND VPWR VPWR _734__786/HI U$$2472/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_94_0 _692__912/HI U$$2190/X U$$2323/X VGND VGND VPWR VPWR dadda_fa_2_95_5/B
+ dadda_fa_2_94_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_150_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$340 final_adder.U$$340/A final_adder.U$$340/B VGND VGND VPWR VPWR
+ final_adder.U$$362/B sky130_fd_sc_hd__and2_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_612_ _612_/CLK _612_/D VGND VGND VPWR VPWR _612_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$362 final_adder.U$$362/A final_adder.U$$362/B VGND VGND VPWR VPWR
+ final_adder.U$$372/A sky130_fd_sc_hd__and2_1
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$201 U$$64/A1 U$$141/X U$$66/A1 U$$142/X VGND VGND VPWR VPWR U$$202/A sky130_fd_sc_hd__a22o_1
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_106_0 dadda_fa_6_106_0/A dadda_fa_6_106_0/B dadda_fa_6_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_107_0/B dadda_fa_7_106_0/CIN sky130_fd_sc_hd__fa_2
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$373 final_adder.U$$372/A final_adder.U$$361/X final_adder.U$$363/X
+ VGND VGND VPWR VPWR final_adder.U$$373/X sky130_fd_sc_hd__a21o_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$212 U$$212/A U$$262/B VGND VGND VPWR VPWR U$$212/X sky130_fd_sc_hd__xor2_2
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$223 U$$86/A1 U$$141/X U$$88/A1 U$$142/X VGND VGND VPWR VPWR U$$224/A sky130_fd_sc_hd__a22o_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$395 final_adder.U$$358/B final_adder.U$$670/B final_adder.U$$333/X
+ VGND VGND VPWR VPWR final_adder.U$$678/B sky130_fd_sc_hd__a21o_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$234 U$$234/A U$$274/A VGND VGND VPWR VPWR U$$234/X sky130_fd_sc_hd__xor2_1
XFILLER_84_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_543_ _543_/CLK _543_/D VGND VGND VPWR VPWR _543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$245 U$$928/B1 U$$141/X _603_/Q U$$142/X VGND VGND VPWR VPWR U$$246/A sky130_fd_sc_hd__a22o_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$256 U$$256/A U$$262/B VGND VGND VPWR VPWR U$$256/X sky130_fd_sc_hd__xor2_1
XFILLER_72_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_3 dadda_fa_3_26_3/A dadda_fa_3_26_3/B dadda_fa_3_26_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_27_1/B dadda_fa_4_26_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_73_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$267 U$$952/A1 U$$141/X U$$952/B1 U$$142/X VGND VGND VPWR VPWR U$$268/A sky130_fd_sc_hd__a22o_1
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$278 U$$276/Y _620_/Q U$$274/A U$$277/X U$$274/Y VGND VGND VPWR VPWR U$$278/X sky130_fd_sc_hd__a32o_4
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$289 U$$289/A U$$357/B VGND VGND VPWR VPWR U$$289/X sky130_fd_sc_hd__xor2_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_474_ _474_/CLK _474_/D VGND VGND VPWR VPWR _474_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_93_0 dadda_fa_6_93_0/A dadda_fa_6_93_0/B dadda_fa_6_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_94_0/B dadda_fa_7_93_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_139_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$6 U$$6/A1 U$$4/X U$$8/A1 U$$5/X VGND VGND VPWR VPWR U$$7/A sky130_fd_sc_hd__a22o_1
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput309 _199_/Q VGND VGND VPWR VPWR o[31] sky130_fd_sc_hd__buf_2
XFILLER_154_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_683__903 VGND VGND VPWR VPWR _683__903/HI _683__903/LO sky130_fd_sc_hd__conb_1
XFILLER_45_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$790 U$$790/A U$$822/A VGND VGND VPWR VPWR U$$790/X sky130_fd_sc_hd__xor2_1
XFILLER_17_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_6 U$$3492/X U$$3625/X U$$3758/X VGND VGND VPWR VPWR dadda_fa_2_81_2/CIN
+ dadda_fa_2_80_5/B sky130_fd_sc_hd__fa_1
XFILLER_132_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_73_5 U$$3877/X U$$4010/X U$$4143/X VGND VGND VPWR VPWR dadda_fa_2_74_2/A
+ dadda_fa_2_73_5/A sky130_fd_sc_hd__fa_1
XFILLER_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_66_4 U$$4129/X U$$4262/X U$$4395/X VGND VGND VPWR VPWR dadda_fa_2_67_1/CIN
+ dadda_fa_2_66_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_3 U$$2785/X U$$2918/X U$$3051/X VGND VGND VPWR VPWR dadda_fa_2_60_1/B
+ dadda_fa_2_59_4/B sky130_fd_sc_hd__fa_1
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_36_2 dadda_fa_4_36_2/A dadda_fa_4_36_2/B dadda_fa_4_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/CIN dadda_fa_5_36_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_29_1 dadda_fa_4_29_1/A dadda_fa_4_29_1/B dadda_fa_4_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/B dadda_fa_5_29_1/B sky130_fd_sc_hd__fa_2
XFILLER_70_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ _333_/CLK _190_/D VGND VGND VPWR VPWR _190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_ha_0_62_5 U$$2126/X U$$2259/X VGND VGND VPWR VPWR dadda_fa_1_63_7/A dadda_fa_2_62_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_135_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4505 U$$4505/A U$$4505/B VGND VGND VPWR VPWR U$$4505/X sky130_fd_sc_hd__xor2_1
XU$$4516 U$$952/B1 U$$4388/X U$$819/A1 U$$4389/X VGND VGND VPWR VPWR U$$4517/A sky130_fd_sc_hd__a22o_1
XFILLER_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_61_3 U$$1326/X U$$1459/X U$$1592/X VGND VGND VPWR VPWR dadda_fa_1_62_6/CIN
+ dadda_fa_1_61_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_708__928 VGND VGND VPWR VPWR _708__928/HI _708__928/LO sky130_fd_sc_hd__conb_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3804 U$$3804/A U$$3835/A VGND VGND VPWR VPWR U$$3804/X sky130_fd_sc_hd__xor2_1
XU$$19 U$$19/A U$$9/B VGND VGND VPWR VPWR U$$19/X sky130_fd_sc_hd__xor2_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3815 U$$4500/A1 U$$3703/X U$$4502/A1 U$$3704/X VGND VGND VPWR VPWR U$$3816/A sky130_fd_sc_hd__a22o_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3826 U$$3826/A U$$3835/A VGND VGND VPWR VPWR U$$3826/X sky130_fd_sc_hd__xor2_1
XFILLER_131_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3837 _672_/Q VGND VGND VPWR VPWR U$$3839/B sky130_fd_sc_hd__inv_1
XFILLER_131_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$170 final_adder.U$$665/A final_adder.U$$664/A VGND VGND VPWR VPWR
+ final_adder.U$$276/A sky130_fd_sc_hd__and2_1
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$181 final_adder.U$$675/A final_adder.U$$547/B1 final_adder.U$$181/B1
+ VGND VGND VPWR VPWR final_adder.U$$181/X sky130_fd_sc_hd__a21o_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_1 dadda_fa_3_31_1/A dadda_fa_3_31_1/B dadda_fa_3_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_0/CIN dadda_fa_4_31_2/A sky130_fd_sc_hd__fa_2
XU$$3848 U$$4122/A1 U$$3912/A2 _555_/Q U$$3912/B2 VGND VGND VPWR VPWR U$$3849/A sky130_fd_sc_hd__a22o_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3859 U$$3859/A U$$3893/B VGND VGND VPWR VPWR U$$3859/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$192 final_adder.U$$687/A final_adder.U$$686/A VGND VGND VPWR VPWR
+ final_adder.U$$288/B sky130_fd_sc_hd__and2_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_24_0 U$$720/X U$$853/X U$$986/X VGND VGND VPWR VPWR dadda_fa_4_25_0/B
+ dadda_fa_4_24_1/CIN sky130_fd_sc_hd__fa_2
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ _532_/CLK _526_/D VGND VGND VPWR VPWR _526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_457_ _464_/CLK _457_/D VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_388_ _535_/CLK _388_/D VGND VGND VPWR VPWR _388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_90_5 dadda_fa_2_90_5/A dadda_fa_2_90_5/B dadda_fa_2_90_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_2/A dadda_fa_4_90_0/A sky130_fd_sc_hd__fa_2
XFILLER_142_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_83_4 dadda_fa_2_83_4/A dadda_fa_2_83_4/B dadda_fa_2_83_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/CIN dadda_fa_3_83_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_3 dadda_fa_2_76_3/A dadda_fa_2_76_3/B dadda_fa_2_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/B dadda_fa_3_76_3/B sky130_fd_sc_hd__fa_1
XFILLER_141_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_69_2 dadda_fa_2_69_2/A dadda_fa_2_69_2/B dadda_fa_2_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/A dadda_fa_3_69_3/A sky130_fd_sc_hd__fa_1
XFILLER_110_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_46_1 dadda_fa_5_46_1/A dadda_fa_5_46_1/B dadda_fa_5_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/B dadda_fa_7_46_0/A sky130_fd_sc_hd__fa_2
XFILLER_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_39_0 dadda_fa_5_39_0/A dadda_fa_5_39_0/B dadda_fa_5_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/A dadda_fa_6_39_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_120_1 dadda_fa_5_120_1/A dadda_fa_5_120_1/B dadda_ha_4_120_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_121_0/B dadda_fa_7_120_0/A sky130_fd_sc_hd__fa_2
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_113_0 dadda_fa_5_113_0/A dadda_fa_5_113_0/B dadda_fa_5_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/A dadda_fa_6_113_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_71_2 U$$2942/X U$$3075/X U$$3208/X VGND VGND VPWR VPWR dadda_fa_2_72_1/A
+ dadda_fa_2_71_4/A sky130_fd_sc_hd__fa_1
XFILLER_8_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_64_1 U$$2928/X U$$3061/X U$$3194/X VGND VGND VPWR VPWR dadda_fa_2_65_0/CIN
+ dadda_fa_2_64_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_41_0 dadda_fa_4_41_0/A dadda_fa_4_41_0/B dadda_fa_4_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/A dadda_fa_5_41_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_57_0 U$$1185/X U$$1318/X U$$1451/X VGND VGND VPWR VPWR dadda_fa_2_58_0/B
+ dadda_fa_2_57_3/B sky130_fd_sc_hd__fa_1
X_846__898 VGND VGND VPWR VPWR _846__898/HI U$$965/A1 sky130_fd_sc_hd__conb_1
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1709 U$$1709/A U$$1739/B VGND VGND VPWR VPWR U$$1709/X sky130_fd_sc_hd__xor2_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _463_/CLK _311_/D VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_242_ _501_/CLK _242_/D VGND VGND VPWR VPWR _242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_173_ _333_/CLK _173_/D VGND VGND VPWR VPWR _173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 a[26] VGND VGND VPWR VPWR _642_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_156_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_93_3 dadda_fa_3_93_3/A dadda_fa_3_93_3/B dadda_fa_3_93_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/B dadda_fa_4_93_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_86_2 dadda_fa_3_86_2/A dadda_fa_3_86_2/B dadda_fa_3_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/A dadda_fa_4_86_2/B sky130_fd_sc_hd__fa_2
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_79_1 dadda_fa_3_79_1/A dadda_fa_3_79_1/B dadda_fa_3_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/CIN dadda_fa_4_79_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_56_0 dadda_fa_6_56_0/A dadda_fa_6_56_0/B dadda_fa_6_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_57_0/B dadda_fa_7_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater609 U$$3/A VGND VGND VPWR VPWR U$$9/B sky130_fd_sc_hd__buf_12
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4302 U$$4302/A U$$4332/B VGND VGND VPWR VPWR U$$4302/X sky130_fd_sc_hd__xor2_1
XU$$4313 _581_/Q U$$4381/A2 _582_/Q U$$4381/B2 VGND VGND VPWR VPWR U$$4314/A sky130_fd_sc_hd__a22o_1
XFILLER_78_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4324 U$$4324/A U$$4384/A VGND VGND VPWR VPWR U$$4324/X sky130_fd_sc_hd__xor2_1
XU$$4335 U$$4335/A1 U$$4377/A2 U$$90/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4336/A sky130_fd_sc_hd__a22o_1
XU$$4346 U$$4346/A _679_/Q VGND VGND VPWR VPWR U$$4346/X sky130_fd_sc_hd__xor2_1
XU$$3601 U$$3601/A U$$3625/B VGND VGND VPWR VPWR U$$3601/X sky130_fd_sc_hd__xor2_1
XFILLER_19_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3612 _573_/Q U$$3668/A2 _574_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3613/A sky130_fd_sc_hd__a22o_1
XU$$4357 U$$4494/A1 U$$4377/A2 U$$4496/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4358/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4368 U$$4368/A U$$4384/A VGND VGND VPWR VPWR U$$4368/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_2 dadda_fa_4_115_2/A dadda_fa_4_115_2/B dadda_fa_4_115_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_116_0/CIN dadda_fa_5_115_1/CIN sky130_fd_sc_hd__fa_1
XU$$3623 U$$3623/A U$$3625/B VGND VGND VPWR VPWR U$$3623/X sky130_fd_sc_hd__xor2_1
XU$$4379 U$$4379/A1 U$$4381/A2 U$$819/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4380/A
+ sky130_fd_sc_hd__a22o_1
XU$$3634 U$$70/B1 U$$3678/A2 U$$759/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3635/A sky130_fd_sc_hd__a22o_1
XU$$2900 U$$2900/A U$$2960/B VGND VGND VPWR VPWR U$$2900/X sky130_fd_sc_hd__xor2_1
XU$$3645 U$$3645/A U$$3699/A VGND VGND VPWR VPWR U$$3645/X sky130_fd_sc_hd__xor2_1
XU$$3656 _595_/Q U$$3668/A2 _596_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3657/A sky130_fd_sc_hd__a22o_1
XU$$2911 U$$3457/B1 U$$2975/A2 U$$4283/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2912/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_108_1 dadda_fa_4_108_1/A dadda_fa_4_108_1/B dadda_fa_4_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/B dadda_fa_5_108_1/B sky130_fd_sc_hd__fa_1
XU$$2922 U$$2922/A U$$2960/B VGND VGND VPWR VPWR U$$2922/X sky130_fd_sc_hd__xor2_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3667 U$$3667/A U$$3699/A VGND VGND VPWR VPWR U$$3667/X sky130_fd_sc_hd__xor2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3678 _606_/Q U$$3678/A2 U$$940/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3679/A sky130_fd_sc_hd__a22o_1
XU$$2933 U$$4303/A1 U$$3009/A2 U$$58/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2934/A sky130_fd_sc_hd__a22o_1
XU$$2944 U$$2944/A U$$3004/B VGND VGND VPWR VPWR U$$2944/X sky130_fd_sc_hd__xor2_1
XU$$3689 U$$3689/A U$$3698/A VGND VGND VPWR VPWR U$$3689/X sky130_fd_sc_hd__xor2_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2955 _587_/Q U$$2881/X _588_/Q U$$2882/X VGND VGND VPWR VPWR U$$2956/A sky130_fd_sc_hd__a22o_1
XFILLER_73_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2966 U$$2966/A U$$3004/B VGND VGND VPWR VPWR U$$2966/X sky130_fd_sc_hd__xor2_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2977 U$$4484/A1 U$$2881/X _599_/Q U$$2882/X VGND VGND VPWR VPWR U$$2978/A sky130_fd_sc_hd__a22o_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2988 U$$2988/A _659_/Q VGND VGND VPWR VPWR U$$2988/X sky130_fd_sc_hd__xor2_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_509_ _509_/CLK _509_/D VGND VGND VPWR VPWR _509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2999 U$$4506/A1 U$$2881/X U$$4508/A1 U$$2882/X VGND VGND VPWR VPWR U$$3000/A sky130_fd_sc_hd__a22o_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_81_1 dadda_fa_2_81_1/A dadda_fa_2_81_1/B dadda_fa_2_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_0/CIN dadda_fa_3_81_2/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_74_0 dadda_fa_2_74_0/A dadda_fa_2_74_0/B dadda_fa_2_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/B dadda_fa_3_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_170_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_50_7 U$$2900/X U$$3033/X U$$3166/X VGND VGND VPWR VPWR dadda_fa_2_51_2/CIN
+ dadda_fa_2_50_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_96_1 dadda_fa_4_96_1/A dadda_fa_4_96_1/B dadda_fa_4_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/B dadda_fa_5_96_1/B sky130_fd_sc_hd__fa_1
XFILLER_137_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_73_0 dadda_fa_7_73_0/A dadda_fa_7_73_0/B dadda_fa_7_73_0/CIN VGND VGND
+ VPWR VPWR _498_/D _369_/D sky130_fd_sc_hd__fa_2
XFILLER_156_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_89_0 dadda_fa_4_89_0/A dadda_fa_4_89_0/B dadda_fa_4_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/A dadda_fa_5_89_1/A sky130_fd_sc_hd__fa_1
XFILLER_152_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2207 U$$2207/A U$$2257/B VGND VGND VPWR VPWR U$$2207/X sky130_fd_sc_hd__xor2_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2218 U$$26/A1 U$$2270/A2 U$$987/A1 U$$2286/B2 VGND VGND VPWR VPWR U$$2219/A sky130_fd_sc_hd__a22o_1
XU$$2229 U$$2229/A U$$2289/B VGND VGND VPWR VPWR U$$2229/X sky130_fd_sc_hd__xor2_1
XU$$1506 _637_/Q VGND VGND VPWR VPWR U$$1506/Y sky130_fd_sc_hd__inv_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1517 U$$8/B1 U$$1591/A2 U$$12/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1518/A sky130_fd_sc_hd__a22o_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1528 U$$1528/A U$$1614/B VGND VGND VPWR VPWR U$$1528/X sky130_fd_sc_hd__xor2_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1539 U$$30/B1 U$$1591/A2 U$$3457/B1 U$$1591/B2 VGND VGND VPWR VPWR U$$1540/A sky130_fd_sc_hd__a22o_1
XFILLER_31_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_225_ _474_/CLK _225_/D VGND VGND VPWR VPWR _225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_91_0 dadda_fa_3_91_0/A dadda_fa_3_91_0/B dadda_fa_3_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/B dadda_fa_4_91_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater406 U$$3668/A2 VGND VGND VPWR VPWR U$$3678/A2 sky130_fd_sc_hd__buf_12
Xrepeater417 U$$2881/X VGND VGND VPWR VPWR U$$3009/A2 sky130_fd_sc_hd__buf_12
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4110 _675_/Q VGND VGND VPWR VPWR U$$4110/Y sky130_fd_sc_hd__inv_1
Xrepeater428 U$$2316/A2 VGND VGND VPWR VPWR U$$2270/A2 sky130_fd_sc_hd__buf_12
Xdadda_fa_2_53_5 dadda_fa_2_53_5/A dadda_fa_2_53_5/B dadda_fa_2_53_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_2/A dadda_fa_4_53_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_120_0 _702__922/HI U$$3971/X U$$4104/X VGND VGND VPWR VPWR dadda_fa_5_121_1/A
+ dadda_fa_5_120_1/B sky130_fd_sc_hd__fa_1
Xrepeater439 U$$1785/X VGND VGND VPWR VPWR U$$1867/A2 sky130_fd_sc_hd__buf_12
XFILLER_93_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4121 U$$4121/A U$$4197/B VGND VGND VPWR VPWR U$$4121/X sky130_fd_sc_hd__xor2_1
XU$$4132 _559_/Q U$$4198/A2 U$$4271/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4133/A sky130_fd_sc_hd__a22o_1
XU$$4143 U$$4143/A U$$4247/A VGND VGND VPWR VPWR U$$4143/X sky130_fd_sc_hd__xor2_1
XU$$4154 U$$4289/B1 U$$4198/A2 U$$4291/B1 U$$4198/B2 VGND VGND VPWR VPWR U$$4155/A
+ sky130_fd_sc_hd__a22o_1
XU$$3420 U$$4379/A1 U$$3292/X U$$819/A1 U$$3293/X VGND VGND VPWR VPWR U$$3421/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_4 dadda_fa_2_46_4/A dadda_fa_2_46_4/B dadda_fa_2_46_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/CIN dadda_fa_3_46_3/CIN sky130_fd_sc_hd__fa_2
XU$$4165 U$$4165/A U$$4247/A VGND VGND VPWR VPWR U$$4165/X sky130_fd_sc_hd__xor2_1
XU$$3431 U$$3431/A1 U$$3429/X U$$8/A1 U$$3430/X VGND VGND VPWR VPWR U$$3432/A sky130_fd_sc_hd__a22o_1
XFILLER_65_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4176 _581_/Q U$$4198/A2 _582_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4177/A sky130_fd_sc_hd__a22o_1
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3442 U$$3442/A U$$3561/A VGND VGND VPWR VPWR U$$3442/X sky130_fd_sc_hd__xor2_1
XFILLER_81_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4187 U$$4187/A U$$4247/A VGND VGND VPWR VPWR U$$4187/X sky130_fd_sc_hd__xor2_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4198 U$$771/B1 U$$4198/A2 U$$912/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4199/A sky130_fd_sc_hd__a22o_1
XU$$3453 _562_/Q U$$3525/A2 _563_/Q U$$3525/B2 VGND VGND VPWR VPWR U$$3454/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_3 U$$2346/X U$$2479/X U$$2612/X VGND VGND VPWR VPWR dadda_fa_3_40_1/B
+ dadda_fa_3_39_3/B sky130_fd_sc_hd__fa_1
XU$$3464 U$$3464/A _667_/Q VGND VGND VPWR VPWR U$$3464/X sky130_fd_sc_hd__xor2_1
XU$$3475 _573_/Q U$$3525/A2 U$$50/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3476/A sky130_fd_sc_hd__a22o_1
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2730 U$$2730/A _655_/Q VGND VGND VPWR VPWR U$$2730/X sky130_fd_sc_hd__xor2_1
XFILLER_74_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2741 _656_/Q VGND VGND VPWR VPWR U$$2743/B sky130_fd_sc_hd__inv_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3486 U$$3486/A U$$3496/B VGND VGND VPWR VPWR U$$3486/X sky130_fd_sc_hd__xor2_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3497 _584_/Q U$$3545/A2 _585_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3498/A sky130_fd_sc_hd__a22o_1
XU$$2752 U$$971/A1 U$$2796/A2 U$$12/B1 U$$2745/X VGND VGND VPWR VPWR U$$2753/A sky130_fd_sc_hd__a22o_1
XU$$2763 U$$2763/A U$$2797/B VGND VGND VPWR VPWR U$$2763/X sky130_fd_sc_hd__xor2_1
XU$$2774 _565_/Q U$$2796/A2 U$$4283/A1 U$$2834/B2 VGND VGND VPWR VPWR U$$2775/A sky130_fd_sc_hd__a22o_1
XU$$2785 U$$2785/A U$$2839/B VGND VGND VPWR VPWR U$$2785/X sky130_fd_sc_hd__xor2_1
XFILLER_34_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2796 U$$56/A1 U$$2796/A2 U$$58/A1 U$$2745/X VGND VGND VPWR VPWR U$$2797/A sky130_fd_sc_hd__a22o_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput209 c[57] VGND VGND VPWR VPWR input209/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$703 final_adder.U$$703/A final_adder.U$$703/B VGND VGND VPWR VPWR
+ _249_/D sky130_fd_sc_hd__xor2_1
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$714 final_adder.U$$714/A final_adder.U$$714/B VGND VGND VPWR VPWR
+ _260_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$725 final_adder.U$$725/A final_adder.U$$725/B VGND VGND VPWR VPWR
+ _271_/D sky130_fd_sc_hd__xor2_1
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$736 final_adder.U$$736/A final_adder.U$$736/B VGND VGND VPWR VPWR
+ _282_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$747 final_adder.U$$747/A final_adder.U$$747/B VGND VGND VPWR VPWR
+ _293_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$608 U$$60/A1 U$$682/A2 U$$62/A1 U$$553/X VGND VGND VPWR VPWR U$$609/A sky130_fd_sc_hd__a22o_1
XU$$619 U$$619/A U$$623/B VGND VGND VPWR VPWR U$$619/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_108_0 U$$3282/X U$$3415/X U$$3548/X VGND VGND VPWR VPWR dadda_fa_4_109_0/B
+ dadda_fa_4_108_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_134_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_56_3 dadda_fa_3_56_3/A dadda_fa_3_56_3/B dadda_fa_3_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/B dadda_fa_4_56_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_49_2 dadda_fa_3_49_2/A dadda_fa_3_49_2/B dadda_fa_3_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/A dadda_fa_4_49_2/B sky130_fd_sc_hd__fa_1
XFILLER_130_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2004 U$$86/A1 U$$2048/A2 U$$88/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$2005/A sky130_fd_sc_hd__a22o_1
XFILLER_114_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2015 U$$2015/A U$$2023/B VGND VGND VPWR VPWR U$$2015/X sky130_fd_sc_hd__xor2_1
XFILLER_74_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_19_0 dadda_fa_6_19_0/A dadda_fa_6_19_0/B dadda_fa_6_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_20_0/B dadda_fa_7_19_0/CIN sky130_fd_sc_hd__fa_1
XU$$2026 U$$930/A1 U$$2052/A2 U$$932/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2027/A sky130_fd_sc_hd__a22o_1
XU$$2037 U$$2037/A U$$2055/A VGND VGND VPWR VPWR U$$2037/X sky130_fd_sc_hd__xor2_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1303 U$$70/A1 U$$1237/X U$$70/B1 U$$1238/X VGND VGND VPWR VPWR U$$1304/A sky130_fd_sc_hd__a22o_1
XU$$2048 U$$4514/A1 U$$2048/A2 _614_/Q U$$2048/B2 VGND VGND VPWR VPWR U$$2049/A sky130_fd_sc_hd__a22o_1
XU$$1314 U$$1314/A U$$1369/A VGND VGND VPWR VPWR U$$1314/X sky130_fd_sc_hd__xor2_1
XU$$2059 U$$2057/Y _646_/Q U$$2055/A U$$2058/X U$$2055/Y VGND VGND VPWR VPWR U$$2059/X
+ sky130_fd_sc_hd__a32o_4
XU$$1325 U$$92/A1 U$$1341/A2 U$$92/B1 U$$1341/B2 VGND VGND VPWR VPWR U$$1326/A sky130_fd_sc_hd__a22o_1
XFILLER_188_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1336 U$$1336/A U$$1336/B VGND VGND VPWR VPWR U$$1336/X sky130_fd_sc_hd__xor2_1
XU$$1347 U$$936/A1 U$$1367/A2 _606_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1348/A sky130_fd_sc_hd__a22o_1
XFILLER_188_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1358 U$$1358/A U$$1369/A VGND VGND VPWR VPWR U$$1358/X sky130_fd_sc_hd__xor2_1
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1369 U$$1369/A VGND VGND VPWR VPWR U$$1369/Y sky130_fd_sc_hd__inv_1
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_208_ _329_/CLK _208_/D VGND VGND VPWR VPWR _208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_51_2 dadda_fa_2_51_2/A dadda_fa_2_51_2/B dadda_fa_2_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/A dadda_fa_3_51_3/A sky130_fd_sc_hd__fa_2
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_44_1 U$$2755/X U$$2888/X U$$3021/X VGND VGND VPWR VPWR dadda_fa_3_45_0/CIN
+ dadda_fa_3_44_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$10 _434_/Q _306_/Q VGND VGND VPWR VPWR final_adder.U$$505/B1 final_adder.U$$632/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$21 _445_/Q _317_/Q VGND VGND VPWR VPWR final_adder.U$$149/B1 final_adder.U$$643/A
+ sky130_fd_sc_hd__ha_1
XU$$3250 U$$3250/A U$$3270/B VGND VGND VPWR VPWR U$$3250/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_21_0 dadda_fa_5_21_0/A dadda_fa_5_21_0/B dadda_fa_5_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/A dadda_fa_6_21_0/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$32 _456_/Q _328_/Q VGND VGND VPWR VPWR final_adder.U$$527/B1 final_adder.U$$654/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_0 U$$746/X U$$879/X U$$1012/X VGND VGND VPWR VPWR dadda_fa_3_38_0/B
+ dadda_fa_3_37_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$43 _467_/Q _339_/Q VGND VGND VPWR VPWR final_adder.U$$171/B1 final_adder.U$$665/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3261 U$$4494/A1 U$$3155/X U$$934/A1 U$$3156/X VGND VGND VPWR VPWR U$$3262/A sky130_fd_sc_hd__a22o_1
XU$$3272 U$$3272/A _663_/Q VGND VGND VPWR VPWR U$$3272/X sky130_fd_sc_hd__xor2_1
XFILLER_81_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$54 _478_/Q _350_/Q VGND VGND VPWR VPWR final_adder.U$$549/B1 final_adder.U$$676/A
+ sky130_fd_sc_hd__ha_1
XU$$3283 U$$4379/A1 U$$3155/X U$$819/A1 U$$3156/X VGND VGND VPWR VPWR U$$3284/A sky130_fd_sc_hd__a22o_1
XFILLER_179_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$65 _489_/Q _361_/Q VGND VGND VPWR VPWR final_adder.U$$193/B1 final_adder.U$$687/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3294 U$$3294/A1 U$$3412/A2 U$$4255/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3295/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$76 _500_/Q _372_/Q VGND VGND VPWR VPWR final_adder.U$$571/B1 final_adder.U$$698/A
+ sky130_fd_sc_hd__ha_1
XFILLER_179_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2560 U$$94/A1 U$$2574/A2 U$$94/B1 U$$2584/B2 VGND VGND VPWR VPWR U$$2561/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$87 _511_/Q _383_/Q VGND VGND VPWR VPWR final_adder.U$$215/B1 final_adder.U$$709/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$98 _522_/Q _394_/Q VGND VGND VPWR VPWR final_adder.U$$593/B1 final_adder.U$$720/A
+ sky130_fd_sc_hd__ha_1
XU$$2571 U$$2571/A U$$2603/A VGND VGND VPWR VPWR U$$2571/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2582 _606_/Q U$$2470/X U$$940/A1 U$$2471/X VGND VGND VPWR VPWR U$$2583/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2593 U$$2593/A U$$2603/A VGND VGND VPWR VPWR U$$2593/X sky130_fd_sc_hd__xor2_1
XFILLER_34_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1870 U$$1870/A U$$1872/B VGND VGND VPWR VPWR U$$1870/X sky130_fd_sc_hd__xor2_1
XU$$1881 _598_/Q U$$1903/A2 _599_/Q U$$1903/B2 VGND VGND VPWR VPWR U$$1882/A sky130_fd_sc_hd__a22o_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1892 U$$1892/A U$$1904/B VGND VGND VPWR VPWR U$$1892/X sky130_fd_sc_hd__xor2_1
XFILLER_30_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_89_3 U$$2978/X U$$3111/X U$$3244/X VGND VGND VPWR VPWR dadda_fa_2_90_4/CIN
+ dadda_fa_3_89_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_66_2 dadda_fa_4_66_2/A dadda_fa_4_66_2/B dadda_fa_4_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/CIN dadda_fa_5_66_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_59_1 dadda_fa_4_59_1/A dadda_fa_4_59_1/B dadda_fa_4_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/B dadda_fa_5_59_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$511 final_adder.U$$638/A final_adder.U$$638/B final_adder.U$$511/B1
+ VGND VGND VPWR VPWR final_adder.U$$639/B sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_36_0 dadda_fa_7_36_0/A dadda_fa_7_36_0/B dadda_fa_7_36_0/CIN VGND VGND
+ VPWR VPWR _461_/D _332_/D sky130_fd_sc_hd__fa_2
XFILLER_69_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$533 final_adder.U$$660/A final_adder.U$$660/B final_adder.U$$533/B1
+ VGND VGND VPWR VPWR final_adder.U$$661/B sky130_fd_sc_hd__a21o_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$555 final_adder.U$$682/A final_adder.U$$682/B final_adder.U$$555/B1
+ VGND VGND VPWR VPWR final_adder.U$$683/B sky130_fd_sc_hd__a21o_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$405 U$$405/A _621_/Q VGND VGND VPWR VPWR U$$405/X sky130_fd_sc_hd__xor2_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$577 final_adder.U$$704/A final_adder.U$$704/B final_adder.U$$577/B1
+ VGND VGND VPWR VPWR final_adder.U$$705/B sky130_fd_sc_hd__a21o_1
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$416 U$$414/B _621_/Q _622_/Q U$$411/Y VGND VGND VPWR VPWR U$$416/X sky130_fd_sc_hd__a22o_4
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$427 U$$16/A1 U$$545/A2 U$$975/B1 U$$416/X VGND VGND VPWR VPWR U$$428/A sky130_fd_sc_hd__a22o_1
XFILLER_84_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$599 final_adder.U$$726/A final_adder.U$$726/B final_adder.U$$599/B1
+ VGND VGND VPWR VPWR final_adder.U$$727/B sky130_fd_sc_hd__a21o_1
XU$$438 U$$438/A U$$530/B VGND VGND VPWR VPWR U$$438/X sky130_fd_sc_hd__xor2_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$449 U$$38/A1 U$$491/A2 U$$40/A1 U$$416/X VGND VGND VPWR VPWR U$$450/A sky130_fd_sc_hd__a22o_1
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_490_ _490_/CLK _490_/D VGND VGND VPWR VPWR _490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_61_1 dadda_fa_3_61_1/A dadda_fa_3_61_1/B dadda_fa_3_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/CIN dadda_fa_4_61_2/A sky130_fd_sc_hd__fa_1
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_0 dadda_fa_3_54_0/A dadda_fa_3_54_0/B dadda_fa_3_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/B dadda_fa_4_54_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$950 U$$950/A1 U$$826/X U$$952/A1 U$$827/X VGND VGND VPWR VPWR U$$951/A sky130_fd_sc_hd__a22o_1
XU$$1100 U$$1098/Y _632_/Q U$$998/B U$$1099/X U$$1096/Y VGND VGND VPWR VPWR U$$1100/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$961 U$$998/B VGND VGND VPWR VPWR U$$961/Y sky130_fd_sc_hd__inv_1
XU$$972 U$$972/A U$$998/B VGND VGND VPWR VPWR U$$972/X sky130_fd_sc_hd__xor2_2
XU$$1111 U$$1111/A U$$1189/B VGND VGND VPWR VPWR U$$1111/X sky130_fd_sc_hd__xor2_1
XFILLER_189_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$983 U$$983/A1 U$$999/A2 U$$26/A1 U$$999/B2 VGND VGND VPWR VPWR U$$984/A sky130_fd_sc_hd__a22o_1
XU$$1122 U$$26/A1 U$$1200/A2 U$$987/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1123/A sky130_fd_sc_hd__a22o_1
XU$$994 U$$994/A U$$998/B VGND VGND VPWR VPWR U$$994/X sky130_fd_sc_hd__xor2_1
XU$$1133 U$$1133/A U$$1189/B VGND VGND VPWR VPWR U$$1133/X sky130_fd_sc_hd__xor2_1
XFILLER_90_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1144 U$$48/A1 U$$1200/A2 U$$50/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1145/A sky130_fd_sc_hd__a22o_1
XU$$1155 U$$1155/A U$$1167/B VGND VGND VPWR VPWR U$$1155/X sky130_fd_sc_hd__xor2_1
XU$$1166 U$$68/B1 U$$1218/A2 U$$72/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1167/A sky130_fd_sc_hd__a22o_1
XU$$1177 U$$1177/A U$$1232/A VGND VGND VPWR VPWR U$$1177/X sky130_fd_sc_hd__xor2_2
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1188 U$$92/A1 U$$1200/A2 U$$94/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1189/A sky130_fd_sc_hd__a22o_1
XU$$1199 U$$1199/A _633_/Q VGND VGND VPWR VPWR U$$1199/X sky130_fd_sc_hd__xor2_1
XFILLER_188_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_111_0 dadda_fa_7_111_0/A dadda_fa_7_111_0/B dadda_fa_7_111_0/CIN VGND
+ VGND VPWR VPWR _536_/D _407_/D sky130_fd_sc_hd__fa_2
XFILLER_15_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_99_2 U$$3264/X U$$3397/X U$$3530/X VGND VGND VPWR VPWR dadda_fa_3_100_1/CIN
+ dadda_fa_3_99_3/B sky130_fd_sc_hd__fa_1
XFILLER_172_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_76_1 dadda_fa_5_76_1/A dadda_fa_5_76_1/B dadda_fa_5_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/B dadda_fa_7_76_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_5_69_0 dadda_fa_5_69_0/A dadda_fa_5_69_0/B dadda_fa_5_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/A dadda_fa_6_69_0/CIN sky130_fd_sc_hd__fa_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_8 dadda_fa_1_68_8/A dadda_fa_1_68_8/B dadda_fa_1_68_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_3/A dadda_fa_3_68_0/A sky130_fd_sc_hd__fa_2
XFILLER_140_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3080 _581_/Q U$$3018/X U$$4178/A1 U$$3019/X VGND VGND VPWR VPWR U$$3081/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_8_0 dadda_fa_6_8_0/A dadda_fa_6_8_0/B dadda_fa_6_8_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_9_0/B dadda_fa_7_8_0/CIN sky130_fd_sc_hd__fa_2
XU$$3091 U$$3091/A U$$3129/B VGND VGND VPWR VPWR U$$3091/X sky130_fd_sc_hd__xor2_1
XU$$2390 U$$2390/A U$$2432/B VGND VGND VPWR VPWR U$$2390/X sky130_fd_sc_hd__xor2_1
XFILLER_167_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_71_0 dadda_fa_4_71_0/A dadda_fa_4_71_0/B dadda_fa_4_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/A dadda_fa_5_71_1/A sky130_fd_sc_hd__fa_1
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_87_0 U$$1643/Y U$$1777/X U$$1910/X VGND VGND VPWR VPWR dadda_fa_2_88_3/A
+ dadda_fa_2_87_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$330 final_adder.U$$330/A final_adder.U$$330/B VGND VGND VPWR VPWR
+ final_adder.U$$356/A sky130_fd_sc_hd__and2_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$341 final_adder.U$$340/A final_adder.U$$297/X final_adder.U$$299/X
+ VGND VGND VPWR VPWR final_adder.U$$341/X sky130_fd_sc_hd__a21o_1
X_611_ _611_/CLK _611_/D VGND VGND VPWR VPWR _611_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$363 final_adder.U$$362/A final_adder.U$$341/X final_adder.U$$343/X
+ VGND VGND VPWR VPWR final_adder.U$$363/X sky130_fd_sc_hd__a21o_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$202 U$$202/A U$$262/B VGND VGND VPWR VPWR U$$202/X sky130_fd_sc_hd__xor2_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$213 U$$759/B1 U$$141/X U$$78/A1 U$$142/X VGND VGND VPWR VPWR U$$214/A sky130_fd_sc_hd__a22o_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$385 final_adder.U$$370/B final_adder.U$$654/B final_adder.U$$357/X
+ VGND VGND VPWR VPWR final_adder.U$$670/B sky130_fd_sc_hd__a21o_4
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$224 U$$224/A U$$262/B VGND VGND VPWR VPWR U$$224/X sky130_fd_sc_hd__xor2_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_542_ _615_/CLK _542_/D VGND VGND VPWR VPWR _542_/Q sky130_fd_sc_hd__dfxtp_1
XU$$235 U$$98/A1 U$$141/X U$$98/B1 U$$142/X VGND VGND VPWR VPWR U$$236/A sky130_fd_sc_hd__a22o_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$246 U$$246/A U$$262/B VGND VGND VPWR VPWR U$$246/X sky130_fd_sc_hd__xor2_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$257 U$$942/A1 U$$141/X U$$944/A1 U$$142/X VGND VGND VPWR VPWR U$$258/A sky130_fd_sc_hd__a22o_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$268 U$$268/A _619_/Q VGND VGND VPWR VPWR U$$268/X sky130_fd_sc_hd__xor2_1
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$279 U$$277/B U$$274/A _620_/Q U$$274/Y VGND VGND VPWR VPWR U$$279/X sky130_fd_sc_hd__a22o_4
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_473_ _480_/CLK _473_/D VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$7 U$$7/A U$$9/B VGND VGND VPWR VPWR U$$7/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_86_0 dadda_fa_6_86_0/A dadda_fa_6_86_0/B dadda_fa_6_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_87_0/B dadda_fa_7_86_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$780 U$$780/A _627_/Q VGND VGND VPWR VPWR U$$780/X sky130_fd_sc_hd__xor2_2
XU$$791 U$$928/A1 U$$817/A2 U$$928/B1 U$$817/B2 VGND VGND VPWR VPWR U$$792/A sky130_fd_sc_hd__a22o_1
XFILLER_90_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR _536_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_192_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_80_7 U$$3891/X U$$4024/X U$$4157/X VGND VGND VPWR VPWR dadda_fa_2_81_3/A
+ dadda_fa_2_80_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_63_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_6 U$$4276/X U$$4409/X input227/X VGND VGND VPWR VPWR dadda_fa_2_74_2/B
+ dadda_fa_2_73_5/B sky130_fd_sc_hd__fa_2
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_66_5 input219/X dadda_fa_1_66_5/B dadda_fa_1_66_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_67_2/A dadda_fa_2_66_5/A sky130_fd_sc_hd__fa_2
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_4 U$$3184/X U$$3317/X U$$3450/X VGND VGND VPWR VPWR dadda_fa_2_60_1/CIN
+ dadda_fa_2_59_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_29_2 dadda_fa_4_29_2/A dadda_fa_4_29_2/B dadda_fa_4_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/CIN dadda_fa_5_29_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_15_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4506 U$$4506/A1 U$$4388/X U$$4508/A1 U$$4389/X VGND VGND VPWR VPWR U$$4507/A sky130_fd_sc_hd__a22o_1
XU$$4517 U$$4517/A U$$4517/B VGND VGND VPWR VPWR U$$4517/X sky130_fd_sc_hd__xor2_2
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3805 U$$654/A1 U$$3703/X U$$4492/A1 U$$3704/X VGND VGND VPWR VPWR U$$3806/A sky130_fd_sc_hd__a22o_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_18_2 U$$841/X U$$974/X VGND VGND VPWR VPWR dadda_fa_4_19_1/CIN dadda_ha_3_18_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3816 U$$3816/A U$$3835/A VGND VGND VPWR VPWR U$$3816/X sky130_fd_sc_hd__xor2_1
XU$$3827 U$$539/A1 U$$3703/X _613_/Q U$$3704/X VGND VGND VPWR VPWR U$$3828/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$160 final_adder.U$$655/A final_adder.U$$654/A VGND VGND VPWR VPWR
+ final_adder.U$$272/B sky130_fd_sc_hd__and2_1
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3838 _673_/Q VGND VGND VPWR VPWR U$$3838/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$171 final_adder.U$$665/A final_adder.U$$537/B1 final_adder.U$$171/B1
+ VGND VGND VPWR VPWR final_adder.U$$171/X sky130_fd_sc_hd__a21o_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3849 U$$3849/A U$$3893/B VGND VGND VPWR VPWR U$$3849/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$182 final_adder.U$$677/A final_adder.U$$676/A VGND VGND VPWR VPWR
+ final_adder.U$$282/A sky130_fd_sc_hd__and2_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_2 dadda_fa_3_31_2/A dadda_fa_3_31_2/B dadda_fa_3_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/A dadda_fa_4_31_2/B sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$193 final_adder.U$$687/A final_adder.U$$559/B1 final_adder.U$$193/B1
+ VGND VGND VPWR VPWR final_adder.U$$193/X sky130_fd_sc_hd__a21o_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_24_1 U$$1119/X U$$1252/X U$$1385/X VGND VGND VPWR VPWR dadda_fa_4_25_0/CIN
+ dadda_fa_4_24_2/A sky130_fd_sc_hd__fa_2
XFILLER_122_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_525_ _537_/CLK _525_/D VGND VGND VPWR VPWR _525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_17_0 U$$41/X U$$174/X U$$307/X VGND VGND VPWR VPWR dadda_fa_4_18_1/B dadda_fa_4_17_2/B
+ sky130_fd_sc_hd__fa_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_456_ _456_/CLK _456_/D VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_387_ _387_/CLK _387_/D VGND VGND VPWR VPWR _387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_83_5 dadda_fa_2_83_5/A dadda_fa_2_83_5/B dadda_fa_2_83_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_2/A dadda_fa_4_83_0/A sky130_fd_sc_hd__fa_2
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_76_4 dadda_fa_2_76_4/A dadda_fa_2_76_4/B dadda_fa_2_76_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/CIN dadda_fa_3_76_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_69_3 dadda_fa_2_69_3/A dadda_fa_2_69_3/B dadda_fa_2_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/B dadda_fa_3_69_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_5_39_1 dadda_fa_5_39_1/A dadda_fa_5_39_1/B dadda_fa_5_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/B dadda_fa_7_39_0/A sky130_fd_sc_hd__fa_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_113_1 dadda_fa_5_113_1/A dadda_fa_5_113_1/B dadda_fa_5_113_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/B dadda_fa_7_113_0/A sky130_fd_sc_hd__fa_1
XFILLER_192_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_106_0 dadda_fa_5_106_0/A dadda_fa_5_106_0/B dadda_fa_5_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/A dadda_fa_6_106_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_71_3 U$$3341/X U$$3474/X U$$3607/X VGND VGND VPWR VPWR dadda_fa_2_72_1/B
+ dadda_fa_2_71_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_64_2 U$$3327/X U$$3460/X U$$3593/X VGND VGND VPWR VPWR dadda_fa_2_65_1/A
+ dadda_fa_2_64_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_41_1 dadda_fa_4_41_1/A dadda_fa_4_41_1/B dadda_fa_4_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/B dadda_fa_5_41_1/B sky130_fd_sc_hd__fa_1
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_1 U$$1584/X U$$1717/X U$$1850/X VGND VGND VPWR VPWR dadda_fa_2_58_0/CIN
+ dadda_fa_2_57_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_28_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_34_0 dadda_fa_4_34_0/A dadda_fa_4_34_0/B dadda_fa_4_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/A dadda_fa_5_34_1/A sky130_fd_sc_hd__fa_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _425_/CLK _310_/D VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_241_ _499_/CLK _241_/D VGND VGND VPWR VPWR _241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_172_ _462_/CLK _172_/D VGND VGND VPWR VPWR _172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_86_3 dadda_fa_3_86_3/A dadda_fa_3_86_3/B dadda_fa_3_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/B dadda_fa_4_86_2/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_79_2 dadda_fa_3_79_2/A dadda_fa_3_79_2/B dadda_fa_3_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/A dadda_fa_4_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_105_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_49_0 dadda_fa_6_49_0/A dadda_fa_6_49_0/B dadda_fa_6_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_50_0/B dadda_fa_7_49_0/CIN sky130_fd_sc_hd__fa_1
XU$$4303 U$$4303/A1 U$$4251/X _577_/Q U$$4252/X VGND VGND VPWR VPWR U$$4304/A sky130_fd_sc_hd__a22o_1
XU$$4314 U$$4314/A _679_/Q VGND VGND VPWR VPWR U$$4314/X sky130_fd_sc_hd__xor2_1
XFILLER_81_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4325 _587_/Q U$$4251/X U$$765/A1 U$$4252/X VGND VGND VPWR VPWR U$$4326/A sky130_fd_sc_hd__a22o_1
XU$$4336 U$$4336/A U$$4384/A VGND VGND VPWR VPWR U$$4336/X sky130_fd_sc_hd__xor2_1
XU$$4347 U$$4484/A1 U$$4377/A2 U$$4486/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4348/A
+ sky130_fd_sc_hd__a22o_1
XU$$3602 U$$4424/A1 U$$3624/A2 U$$4289/A1 U$$3624/B2 VGND VGND VPWR VPWR U$$3603/A
+ sky130_fd_sc_hd__a22o_1
XU$$3613 U$$3613/A U$$3699/A VGND VGND VPWR VPWR U$$3613/X sky130_fd_sc_hd__xor2_1
XU$$4358 U$$4358/A U$$4384/A VGND VGND VPWR VPWR U$$4358/X sky130_fd_sc_hd__xor2_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3624 U$$3624/A1 U$$3624/A2 _580_/Q U$$3624/B2 VGND VGND VPWR VPWR U$$3625/A sky130_fd_sc_hd__a22o_1
XU$$4369 U$$4506/A1 U$$4377/A2 U$$4508/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4370/A
+ sky130_fd_sc_hd__a22o_1
XU$$3635 U$$3635/A _669_/Q VGND VGND VPWR VPWR U$$3635/X sky130_fd_sc_hd__xor2_1
XU$$2901 U$$4271/A1 U$$2975/A2 U$$4273/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2902/A
+ sky130_fd_sc_hd__a22o_1
XU$$3646 _590_/Q U$$3668/A2 _591_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3647/A sky130_fd_sc_hd__a22o_1
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3657 U$$3657/A U$$3699/A VGND VGND VPWR VPWR U$$3657/X sky130_fd_sc_hd__xor2_1
XU$$2912 U$$2912/A U$$2996/B VGND VGND VPWR VPWR U$$2912/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_108_2 dadda_fa_4_108_2/A dadda_fa_4_108_2/B dadda_fa_4_108_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/CIN dadda_fa_5_108_1/CIN sky130_fd_sc_hd__fa_1
XU$$2923 U$$868/A1 U$$3009/A2 U$$48/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2924/A sky130_fd_sc_hd__a22o_1
XU$$3668 _601_/Q U$$3668/A2 U$$928/B1 U$$3668/B2 VGND VGND VPWR VPWR U$$3669/A sky130_fd_sc_hd__a22o_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3679 U$$3679/A _669_/Q VGND VGND VPWR VPWR U$$3679/X sky130_fd_sc_hd__xor2_1
XFILLER_93_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2934 U$$2934/A U$$2996/B VGND VGND VPWR VPWR U$$2934/X sky130_fd_sc_hd__xor2_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2945 U$$4178/A1 U$$2881/X _583_/Q U$$2882/X VGND VGND VPWR VPWR U$$2946/A sky130_fd_sc_hd__a22o_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2956 U$$2956/A U$$3004/B VGND VGND VPWR VPWR U$$2956/X sky130_fd_sc_hd__xor2_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2967 _593_/Q U$$2881/X _594_/Q U$$2882/X VGND VGND VPWR VPWR U$$2968/A sky130_fd_sc_hd__a22o_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2978 U$$2978/A U$$3004/B VGND VGND VPWR VPWR U$$2978/X sky130_fd_sc_hd__xor2_1
XFILLER_178_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_508_ _510_/CLK _508_/D VGND VGND VPWR VPWR _508_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2989 _604_/Q U$$2881/X _605_/Q U$$2882/X VGND VGND VPWR VPWR U$$2990/A sky130_fd_sc_hd__a22o_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ _463_/CLK _439_/D VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _379_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_81_2 dadda_fa_2_81_2/A dadda_fa_2_81_2/B dadda_fa_2_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/A dadda_fa_3_81_3/A sky130_fd_sc_hd__fa_1
XFILLER_138_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_1 dadda_fa_2_74_1/A dadda_fa_2_74_1/B dadda_fa_2_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/CIN dadda_fa_3_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_51_0 dadda_fa_5_51_0/A dadda_fa_5_51_0/B dadda_fa_5_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/A dadda_fa_6_51_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_67_0 dadda_fa_2_67_0/A dadda_fa_2_67_0/B dadda_fa_2_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/B dadda_fa_3_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_clk _369_/CLK VGND VGND VPWR VPWR _488_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_772__824 VGND VGND VPWR VPWR _772__824/HI U$$4390/A1 sky130_fd_sc_hd__conb_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_96_2 dadda_fa_4_96_2/A dadda_fa_4_96_2/B dadda_fa_4_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/CIN dadda_fa_5_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_89_1 dadda_fa_4_89_1/A dadda_fa_4_89_1/B dadda_fa_4_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/B dadda_fa_5_89_1/B sky130_fd_sc_hd__fa_1
X_813__865 VGND VGND VPWR VPWR _813__865/HI U$$4471/B sky130_fd_sc_hd__conb_1
XFILLER_69_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_66_0 dadda_fa_7_66_0/A dadda_fa_7_66_0/B dadda_fa_7_66_0/CIN VGND VGND
+ VPWR VPWR _491_/D _362_/D sky130_fd_sc_hd__fa_2
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2208 U$$16/A1 U$$2196/X U$$18/A1 U$$2197/X VGND VGND VPWR VPWR U$$2209/A sky130_fd_sc_hd__a22o_1
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2219 U$$2219/A U$$2257/B VGND VGND VPWR VPWR U$$2219/X sky130_fd_sc_hd__xor2_1
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1507 _637_/Q VGND VGND VPWR VPWR U$$1507/Y sky130_fd_sc_hd__inv_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1518 U$$1518/A U$$1580/B VGND VGND VPWR VPWR U$$1518/X sky130_fd_sc_hd__xor2_1
XU$$1529 U$$22/A1 U$$1511/X _560_/Q U$$1512/X VGND VGND VPWR VPWR U$$1530/A sky130_fd_sc_hd__a22o_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_22_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _456_/CLK sky130_fd_sc_hd__clkbuf_16
X_224_ _474_/CLK _224_/D VGND VGND VPWR VPWR _224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_91_1 dadda_fa_3_91_1/A dadda_fa_3_91_1/B dadda_fa_3_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/CIN dadda_fa_4_91_2/A sky130_fd_sc_hd__fa_2
XFILLER_100_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_84_0 dadda_fa_3_84_0/A dadda_fa_3_84_0/B dadda_fa_3_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/B dadda_fa_4_84_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_124_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _366_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater407 U$$3566/X VGND VGND VPWR VPWR U$$3668/A2 sky130_fd_sc_hd__buf_12
Xrepeater418 U$$2744/X VGND VGND VPWR VPWR U$$2796/A2 sky130_fd_sc_hd__buf_12
XU$$4100 U$$4100/A U$$4109/A VGND VGND VPWR VPWR U$$4100/X sky130_fd_sc_hd__xor2_1
Xrepeater429 U$$2316/A2 VGND VGND VPWR VPWR U$$2326/A2 sky130_fd_sc_hd__buf_12
XU$$4111 _676_/Q VGND VGND VPWR VPWR U$$4113/B sky130_fd_sc_hd__inv_1
XU$$4122 U$$4122/A1 U$$4198/A2 _555_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4123/A sky130_fd_sc_hd__a22o_1
XU$$4133 U$$4133/A U$$4247/A VGND VGND VPWR VPWR U$$4133/X sky130_fd_sc_hd__xor2_1
XFILLER_66_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4144 _565_/Q U$$4244/A2 _566_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4145/A sky130_fd_sc_hd__a22o_1
XFILLER_168_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3410 U$$4506/A1 U$$3412/A2 U$$4508/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3411/A
+ sky130_fd_sc_hd__a22o_1
XU$$4155 U$$4155/A U$$4247/A VGND VGND VPWR VPWR U$$4155/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_0 U$$4223/X U$$4356/X U$$4489/X VGND VGND VPWR VPWR dadda_fa_5_114_0/A
+ dadda_fa_5_113_1/A sky130_fd_sc_hd__fa_2
XU$$3421 U$$3421/A _665_/Q VGND VGND VPWR VPWR U$$3421/X sky130_fd_sc_hd__xor2_1
XU$$4166 U$$4303/A1 U$$4198/A2 _577_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4167/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_5 dadda_fa_2_46_5/A dadda_fa_2_46_5/B dadda_fa_2_46_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_2/A dadda_fa_4_46_0/A sky130_fd_sc_hd__fa_2
XU$$3432 U$$3432/A U$$3561/A VGND VGND VPWR VPWR U$$3432/X sky130_fd_sc_hd__xor2_1
XU$$4177 U$$4177/A U$$4247/A VGND VGND VPWR VPWR U$$4177/X sky130_fd_sc_hd__xor2_1
XU$$3443 U$$975/B1 U$$3429/X U$$842/A1 U$$3430/X VGND VGND VPWR VPWR U$$3444/A sky130_fd_sc_hd__a22o_1
XU$$4188 _587_/Q U$$4114/X U$$765/A1 U$$4115/X VGND VGND VPWR VPWR U$$4189/A sky130_fd_sc_hd__a22o_1
XFILLER_19_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_39_4 input189/X dadda_fa_2_39_4/B dadda_fa_2_39_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_40_1/CIN dadda_fa_3_39_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4199 U$$4199/A U$$4247/A VGND VGND VPWR VPWR U$$4199/X sky130_fd_sc_hd__xor2_1
XU$$3454 U$$3454/A U$$3496/B VGND VGND VPWR VPWR U$$3454/X sky130_fd_sc_hd__xor2_1
XU$$2720 U$$2720/A _655_/Q VGND VGND VPWR VPWR U$$2720/X sky130_fd_sc_hd__xor2_1
XU$$3465 U$$4424/A1 U$$3545/A2 U$$4289/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3466/A
+ sky130_fd_sc_hd__a22o_1
XU$$3476 U$$3476/A U$$3496/B VGND VGND VPWR VPWR U$$3476/X sky130_fd_sc_hd__xor2_1
XU$$2731 _612_/Q U$$2607/X _613_/Q U$$2608/X VGND VGND VPWR VPWR U$$2732/A sky130_fd_sc_hd__a22o_1
XU$$3487 U$$3624/A1 U$$3545/A2 _580_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3488/A sky130_fd_sc_hd__a22o_1
XU$$2742 _657_/Q VGND VGND VPWR VPWR U$$2742/Y sky130_fd_sc_hd__inv_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3498 U$$3498/A U$$3536/B VGND VGND VPWR VPWR U$$3498/X sky130_fd_sc_hd__xor2_1
XU$$2753 U$$2753/A U$$2797/B VGND VGND VPWR VPWR U$$2753/X sky130_fd_sc_hd__xor2_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2764 U$$983/A1 U$$2796/A2 _561_/Q U$$2826/B2 VGND VGND VPWR VPWR U$$2765/A sky130_fd_sc_hd__a22o_1
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2775 U$$2775/A U$$2839/B VGND VGND VPWR VPWR U$$2775/X sky130_fd_sc_hd__xor2_1
XU$$2786 U$$4291/B1 U$$2870/A2 U$$4156/B1 U$$2834/B2 VGND VGND VPWR VPWR U$$2787/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2797 U$$2797/A U$$2797/B VGND VGND VPWR VPWR U$$2797/X sky130_fd_sc_hd__xor2_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_756__808 VGND VGND VPWR VPWR _756__808/HI U$$3842/A1 sky130_fd_sc_hd__conb_1
XFILLER_57_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _463_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_99_0 dadda_fa_5_99_0/A dadda_fa_5_99_0/B dadda_fa_5_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/A dadda_fa_6_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$704 final_adder.U$$704/A final_adder.U$$704/B VGND VGND VPWR VPWR
+ _250_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$715 final_adder.U$$715/A final_adder.U$$715/B VGND VGND VPWR VPWR
+ _261_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$726 final_adder.U$$726/A final_adder.U$$726/B VGND VGND VPWR VPWR
+ _272_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$737 final_adder.U$$737/A final_adder.U$$737/B VGND VGND VPWR VPWR
+ _283_/D sky130_fd_sc_hd__xor2_1
XFILLER_99_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$748 final_adder.U$$748/A final_adder.U$$748/B VGND VGND VPWR VPWR
+ _294_/D sky130_fd_sc_hd__xor2_2
XFILLER_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$609 U$$609/A U$$661/B VGND VGND VPWR VPWR U$$609/X sky130_fd_sc_hd__xor2_1
XFILLER_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_108_1 U$$3681/X U$$3814/X U$$3947/X VGND VGND VPWR VPWR dadda_fa_4_109_0/CIN
+ dadda_fa_4_108_2/A sky130_fd_sc_hd__fa_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 _182_/Q VGND VGND VPWR VPWR o[14] sky130_fd_sc_hd__buf_2
XFILLER_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_49_3 dadda_fa_3_49_3/A dadda_fa_3_49_3/B dadda_fa_3_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/B dadda_fa_4_49_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2005 U$$2005/A U$$2023/B VGND VGND VPWR VPWR U$$2005/X sky130_fd_sc_hd__xor2_1
XU$$2016 _597_/Q U$$2036/A2 _598_/Q U$$2036/B2 VGND VGND VPWR VPWR U$$2017/A sky130_fd_sc_hd__a22o_1
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2027 U$$2027/A U$$2055/A VGND VGND VPWR VPWR U$$2027/X sky130_fd_sc_hd__xor2_1
XU$$2038 U$$4504/A1 U$$2052/A2 U$$944/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2039/A
+ sky130_fd_sc_hd__a22o_1
XU$$1304 U$$1304/A U$$1336/B VGND VGND VPWR VPWR U$$1304/X sky130_fd_sc_hd__xor2_1
XFILLER_16_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2049 U$$2049/A U$$2055/A VGND VGND VPWR VPWR U$$2049/X sky130_fd_sc_hd__xor2_1
XU$$1315 U$$902/B1 U$$1367/A2 U$$84/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1316/A sky130_fd_sc_hd__a22o_1
XU$$1326 U$$1326/A U$$1342/B VGND VGND VPWR VPWR U$$1326/X sky130_fd_sc_hd__xor2_1
XFILLER_188_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1337 U$$926/A1 U$$1367/A2 _601_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1338/A sky130_fd_sc_hd__a22o_1
XU$$1348 U$$1348/A U$$1369/A VGND VGND VPWR VPWR U$$1348/X sky130_fd_sc_hd__xor2_1
XU$$1359 U$$4510/A1 U$$1367/A2 _612_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1360/A sky130_fd_sc_hd__a22o_1
XFILLER_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_207_ _333_/CLK _207_/D VGND VGND VPWR VPWR _207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_2_clk _431_/CLK VGND VGND VPWR VPWR _438_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_51_3 dadda_fa_2_51_3/A dadda_fa_2_51_3/B dadda_fa_2_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/B dadda_fa_3_51_3/B sky130_fd_sc_hd__fa_2
Xdadda_fa_2_44_2 U$$3129/B input195/X dadda_fa_2_44_2/CIN VGND VGND VPWR VPWR dadda_fa_3_45_1/A
+ dadda_fa_3_44_3/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$11 _435_/Q _307_/Q VGND VGND VPWR VPWR final_adder.U$$139/B1 final_adder.U$$633/A
+ sky130_fd_sc_hd__ha_1
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3240 U$$3240/A _663_/Q VGND VGND VPWR VPWR U$$3240/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_21_1 dadda_fa_5_21_1/A dadda_fa_5_21_1/B dadda_fa_5_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/B dadda_fa_7_21_0/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$22 _446_/Q _318_/Q VGND VGND VPWR VPWR final_adder.U$$517/B1 final_adder.U$$644/A
+ sky130_fd_sc_hd__ha_1
XU$$3251 U$$98/B1 U$$3155/X U$$4486/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3252/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$33 _457_/Q _329_/Q VGND VGND VPWR VPWR final_adder.U$$161/B1 final_adder.U$$655/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3262 U$$3262/A _663_/Q VGND VGND VPWR VPWR U$$3262/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_37_1 U$$1145/X U$$1278/X U$$1411/X VGND VGND VPWR VPWR dadda_fa_3_38_0/CIN
+ dadda_fa_3_37_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$44 _468_/Q _340_/Q VGND VGND VPWR VPWR final_adder.U$$539/B1 final_adder.U$$666/A
+ sky130_fd_sc_hd__ha_1
XU$$3273 U$$4506/A1 U$$3155/X U$$4508/A1 U$$3156/X VGND VGND VPWR VPWR U$$3274/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$55 _479_/Q _351_/Q VGND VGND VPWR VPWR final_adder.U$$183/B1 final_adder.U$$677/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$66 _490_/Q _362_/Q VGND VGND VPWR VPWR final_adder.U$$561/B1 final_adder.U$$688/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3284 U$$3284/A _663_/Q VGND VGND VPWR VPWR U$$3284/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_0 dadda_fa_5_14_0/A dadda_fa_5_14_0/B dadda_fa_5_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/A dadda_fa_6_14_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_81_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2550 _590_/Q U$$2584/A2 U$$908/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2551/A sky130_fd_sc_hd__a22o_1
XU$$3295 U$$3295/A U$$3413/B VGND VGND VPWR VPWR U$$3295/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$77 _501_/Q _373_/Q VGND VGND VPWR VPWR final_adder.U$$205/B1 final_adder.U$$699/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2561 U$$2561/A _653_/Q VGND VGND VPWR VPWR U$$2561/X sky130_fd_sc_hd__xor2_1
XFILLER_179_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$88 _512_/Q _384_/Q VGND VGND VPWR VPWR final_adder.U$$583/B1 final_adder.U$$710/A
+ sky130_fd_sc_hd__ha_2
XU$$2572 _601_/Q U$$2584/A2 U$$928/B1 U$$2584/B2 VGND VGND VPWR VPWR U$$2573/A sky130_fd_sc_hd__a22o_1
XFILLER_110_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$99 _523_/Q _395_/Q VGND VGND VPWR VPWR final_adder.U$$227/B1 final_adder.U$$721/A
+ sky130_fd_sc_hd__ha_2
XFILLER_34_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2583 U$$2583/A _653_/Q VGND VGND VPWR VPWR U$$2583/X sky130_fd_sc_hd__xor2_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2594 U$$950/A1 U$$2470/X U$$4514/A1 U$$2471/X VGND VGND VPWR VPWR U$$2595/A sky130_fd_sc_hd__a22o_1
XU$$1860 U$$1860/A U$$1872/B VGND VGND VPWR VPWR U$$1860/X sky130_fd_sc_hd__xor2_1
XU$$1871 U$$912/A1 U$$1897/A2 U$$914/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1872/A sky130_fd_sc_hd__a22o_1
XU$$1882 U$$1882/A U$$1904/B VGND VGND VPWR VPWR U$$1882/X sky130_fd_sc_hd__xor2_1
XU$$1893 U$$934/A1 U$$1785/X U$$936/A1 U$$1786/X VGND VGND VPWR VPWR U$$1894/A sky130_fd_sc_hd__a22o_1
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_40_3 U$$1284/X U$$1417/X VGND VGND VPWR VPWR dadda_fa_2_41_4/CIN dadda_fa_3_40_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_59_2 dadda_fa_4_59_2/A dadda_fa_4_59_2/B dadda_fa_4_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/CIN dadda_fa_5_59_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$501 final_adder.U$$628/A final_adder.U$$628/B final_adder.U$$6/COUT
+ VGND VGND VPWR VPWR final_adder.U$$629/B sky130_fd_sc_hd__a21o_1
XFILLER_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$523 final_adder.U$$650/A final_adder.U$$650/B final_adder.U$$523/B1
+ VGND VGND VPWR VPWR final_adder.U$$651/B sky130_fd_sc_hd__a21o_1
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_4_10_1 U$$426/X U$$559/X VGND VGND VPWR VPWR dadda_fa_5_11_1/A dadda_ha_4_10_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_85_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$545 final_adder.U$$672/A final_adder.U$$672/B final_adder.U$$545/B1
+ VGND VGND VPWR VPWR final_adder.U$$673/B sky130_fd_sc_hd__a21o_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater760 U$$4255/A1 VGND VGND VPWR VPWR U$$8/A1 sky130_fd_sc_hd__buf_12
Xdadda_fa_7_29_0 dadda_fa_7_29_0/A dadda_fa_7_29_0/B dadda_fa_7_29_0/CIN VGND VGND
+ VPWR VPWR _454_/D _325_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$567 final_adder.U$$694/A final_adder.U$$694/B final_adder.U$$567/B1
+ VGND VGND VPWR VPWR final_adder.U$$695/B sky130_fd_sc_hd__a21o_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$406 U$$952/B1 U$$278/X U$$819/A1 U$$279/X VGND VGND VPWR VPWR U$$407/A sky130_fd_sc_hd__a22o_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$417 U$$417/A1 U$$491/A2 U$$8/A1 U$$416/X VGND VGND VPWR VPWR U$$418/A sky130_fd_sc_hd__a22o_1
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$589 final_adder.U$$716/A final_adder.U$$716/B final_adder.U$$589/B1
+ VGND VGND VPWR VPWR final_adder.U$$717/B sky130_fd_sc_hd__a21o_1
XFILLER_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$428 U$$428/A U$$530/B VGND VGND VPWR VPWR U$$428/X sky130_fd_sc_hd__xor2_1
XFILLER_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$439 U$$987/A1 U$$491/A2 U$$28/B1 U$$416/X VGND VGND VPWR VPWR U$$440/A sky130_fd_sc_hd__a22o_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_778__830 VGND VGND VPWR VPWR _778__830/HI U$$4401/B sky130_fd_sc_hd__conb_1
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_819__871 VGND VGND VPWR VPWR _819__871/HI U$$4483/B sky130_fd_sc_hd__conb_1
XFILLER_138_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_61_2 dadda_fa_3_61_2/A dadda_fa_3_61_2/B dadda_fa_3_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/A dadda_fa_4_61_2/B sky130_fd_sc_hd__fa_1
XFILLER_94_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_1 dadda_fa_3_54_1/A dadda_fa_3_54_1/B dadda_fa_3_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/CIN dadda_fa_4_54_2/A sky130_fd_sc_hd__fa_1
XFILLER_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_31_0 dadda_fa_6_31_0/A dadda_fa_6_31_0/B dadda_fa_6_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_32_0/B dadda_fa_7_31_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_47_0 dadda_fa_3_47_0/A dadda_fa_3_47_0/B dadda_fa_3_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/B dadda_fa_4_47_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_48_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$940 U$$940/A1 U$$826/X U$$942/A1 U$$827/X VGND VGND VPWR VPWR U$$941/A sky130_fd_sc_hd__a22o_1
XU$$951 U$$951/A U$$959/A VGND VGND VPWR VPWR U$$951/X sky130_fd_sc_hd__xor2_1
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$962 U$$998/B U$$962/B VGND VGND VPWR VPWR U$$962/X sky130_fd_sc_hd__and2_1
XU$$1101 U$$1099/B U$$998/B _632_/Q U$$1096/Y VGND VGND VPWR VPWR U$$1101/X sky130_fd_sc_hd__a22o_4
XU$$973 U$$12/B1 U$$999/A2 U$$16/A1 U$$999/B2 VGND VGND VPWR VPWR U$$974/A sky130_fd_sc_hd__a22o_1
XFILLER_91_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1112 U$$14/B1 U$$1200/A2 U$$4265/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1113/A sky130_fd_sc_hd__a22o_1
XU$$1123 U$$1123/A U$$1189/B VGND VGND VPWR VPWR U$$1123/X sky130_fd_sc_hd__xor2_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$984 U$$984/A U$$992/B VGND VGND VPWR VPWR U$$984/X sky130_fd_sc_hd__xor2_1
XFILLER_188_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$995 U$$36/A1 U$$963/X U$$38/A1 U$$999/B2 VGND VGND VPWR VPWR U$$996/A sky130_fd_sc_hd__a22o_1
XU$$1134 U$$38/A1 U$$1200/A2 U$$3191/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1135/A sky130_fd_sc_hd__a22o_1
XFILLER_71_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1145 U$$1145/A U$$1167/B VGND VGND VPWR VPWR U$$1145/X sky130_fd_sc_hd__xor2_1
XU$$1156 U$$60/A1 U$$1200/A2 U$$62/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1157/A sky130_fd_sc_hd__a22o_1
XU$$1167 U$$1167/A U$$1167/B VGND VGND VPWR VPWR U$$1167/X sky130_fd_sc_hd__xor2_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1178 U$$902/B1 U$$1218/A2 U$$84/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1179/A sky130_fd_sc_hd__a22o_1
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1189 U$$1189/A U$$1189/B VGND VGND VPWR VPWR U$$1189/X sky130_fd_sc_hd__xor2_1
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_104_0 dadda_fa_7_104_0/A dadda_fa_7_104_0/B dadda_fa_7_104_0/CIN VGND
+ VGND VPWR VPWR _529_/D _400_/D sky130_fd_sc_hd__fa_2
XFILLER_129_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_3 U$$3663/X U$$3796/X U$$3929/X VGND VGND VPWR VPWR dadda_fa_3_100_2/A
+ dadda_fa_3_99_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_172_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_69_1 dadda_fa_5_69_1/A dadda_fa_5_69_1/B dadda_fa_5_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/B dadda_fa_7_69_0/A sky130_fd_sc_hd__fa_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3070 U$$4303/A1 U$$3090/A2 U$$880/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3071/A
+ sky130_fd_sc_hd__a22o_1
XU$$3081 U$$3081/A U$$3137/B VGND VGND VPWR VPWR U$$3081/X sky130_fd_sc_hd__xor2_1
XU$$3092 U$$76/B1 U$$3146/A2 U$$902/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3093/A sky130_fd_sc_hd__a22o_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2380 U$$2380/A U$$2436/B VGND VGND VPWR VPWR U$$2380/X sky130_fd_sc_hd__xor2_1
XFILLER_50_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2391 U$$4446/A1 U$$2421/A2 U$$3900/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2392/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1690 U$$4291/B1 U$$1726/A2 U$$48/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1691/A sky130_fd_sc_hd__a22o_1
XFILLER_22_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_71_1 dadda_fa_4_71_1/A dadda_fa_4_71_1/B dadda_fa_4_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/B dadda_fa_5_71_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_1 U$$2043/X U$$2176/X U$$2309/X VGND VGND VPWR VPWR dadda_fa_2_88_3/B
+ dadda_fa_2_87_5/A sky130_fd_sc_hd__fa_1
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_64_0 dadda_fa_4_64_0/A dadda_fa_4_64_0/B dadda_fa_4_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/A dadda_fa_5_64_1/A sky130_fd_sc_hd__fa_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_610_ _611_/CLK _610_/D VGND VGND VPWR VPWR _610_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$331 final_adder.U$$330/A final_adder.U$$277/X final_adder.U$$279/X
+ VGND VGND VPWR VPWR final_adder.U$$331/X sky130_fd_sc_hd__a21o_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$342 final_adder.U$$342/A final_adder.U$$342/B VGND VGND VPWR VPWR
+ final_adder.U$$362/A sky130_fd_sc_hd__and2_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$353 final_adder.U$$322/X final_adder.U$$630/B final_adder.U$$323/X
+ VGND VGND VPWR VPWR final_adder.U$$638/B sky130_fd_sc_hd__a21o_2
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$364 final_adder.U$$364/A final_adder.U$$364/B VGND VGND VPWR VPWR
+ final_adder.U$$364/X sky130_fd_sc_hd__and2_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$203 U$$66/A1 U$$141/X U$$68/A1 U$$142/X VGND VGND VPWR VPWR U$$204/A sky130_fd_sc_hd__a22o_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$214 U$$214/A U$$274/A VGND VGND VPWR VPWR U$$214/X sky130_fd_sc_hd__xor2_1
XFILLER_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_541_ _543_/CLK _541_/D VGND VGND VPWR VPWR _541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater590 U$$998/B VGND VGND VPWR VPWR U$$992/B sky130_fd_sc_hd__buf_12
XU$$225 U$$88/A1 U$$141/X U$$90/A1 U$$142/X VGND VGND VPWR VPWR U$$226/A sky130_fd_sc_hd__a22o_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$397 final_adder.U$$360/B final_adder.U$$686/B final_adder.U$$337/X
+ VGND VGND VPWR VPWR final_adder.U$$694/B sky130_fd_sc_hd__a21o_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$236 U$$236/A U$$274/A VGND VGND VPWR VPWR U$$236/X sky130_fd_sc_hd__xor2_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$247 _603_/Q U$$141/X U$$934/A1 U$$142/X VGND VGND VPWR VPWR U$$248/A sky130_fd_sc_hd__a22o_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$258 U$$258/A U$$262/B VGND VGND VPWR VPWR U$$258/X sky130_fd_sc_hd__xor2_1
XU$$269 U$$952/B1 U$$141/X U$$819/A1 U$$142/X VGND VGND VPWR VPWR U$$270/A sky130_fd_sc_hd__a22o_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_472_ _476_/CLK _472_/D VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$8 U$$8/A1 U$$4/X U$$8/B1 U$$5/X VGND VGND VPWR VPWR U$$9/A sky130_fd_sc_hd__a22o_1
XFILLER_154_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_76_1 U$$1223/X U$$1356/X VGND VGND VPWR VPWR dadda_fa_1_77_8/CIN dadda_fa_2_76_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_79_0 dadda_fa_6_79_0/A dadda_fa_6_79_0/B dadda_fa_6_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_80_0/B dadda_fa_7_79_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_141_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$770 U$$770/A U$$778/B VGND VGND VPWR VPWR U$$770/X sky130_fd_sc_hd__xor2_1
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$781 U$$96/A1 U$$785/A2 U$$96/B1 U$$785/B2 VGND VGND VPWR VPWR U$$782/A sky130_fd_sc_hd__a22o_1
XFILLER_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$792 U$$792/A _627_/Q VGND VGND VPWR VPWR U$$792/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_81_0 dadda_fa_5_81_0/A dadda_fa_5_81_0/B dadda_fa_5_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/A dadda_fa_6_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_97_0 U$$2328/Y U$$2462/X U$$2595/X VGND VGND VPWR VPWR dadda_fa_3_98_0/B
+ dadda_fa_3_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_172_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_73_7 dadda_fa_1_73_7/A dadda_fa_1_73_7/B dadda_fa_1_73_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_2/CIN dadda_fa_2_73_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_66_6 dadda_fa_1_66_6/A dadda_fa_1_66_6/B dadda_fa_1_66_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/B dadda_fa_2_66_5/B sky130_fd_sc_hd__fa_1
XFILLER_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_5 U$$3583/X U$$3716/X U$$3849/X VGND VGND VPWR VPWR dadda_fa_2_60_2/A
+ dadda_fa_2_59_5/A sky130_fd_sc_hd__fa_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_740__792 VGND VGND VPWR VPWR _740__792/HI U$$280/A1 sky130_fd_sc_hd__conb_1
XFILLER_167_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_96_0 dadda_fa_7_96_0/A dadda_fa_7_96_0/B dadda_fa_7_96_0/CIN VGND VGND
+ VPWR VPWR _521_/D _392_/D sky130_fd_sc_hd__fa_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4507 U$$4507/A U$$4507/B VGND VGND VPWR VPWR U$$4507/X sky130_fd_sc_hd__xor2_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_111_0 dadda_fa_6_111_0/A dadda_fa_6_111_0/B dadda_fa_6_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_112_0/B dadda_fa_7_111_0/CIN sky130_fd_sc_hd__fa_2
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3806 U$$3806/A U$$3835/A VGND VGND VPWR VPWR U$$3806/X sky130_fd_sc_hd__xor2_1
XFILLER_131_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3817 U$$4502/A1 U$$3703/X U$$4504/A1 U$$3704/X VGND VGND VPWR VPWR U$$3818/A sky130_fd_sc_hd__a22o_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$150 final_adder.U$$645/A final_adder.U$$644/A VGND VGND VPWR VPWR
+ final_adder.U$$266/A sky130_fd_sc_hd__and2_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3828 U$$3828/A U$$3835/A VGND VGND VPWR VPWR U$$3828/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$161 final_adder.U$$655/A final_adder.U$$527/B1 final_adder.U$$161/B1
+ VGND VGND VPWR VPWR final_adder.U$$161/X sky130_fd_sc_hd__a21o_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$172 final_adder.U$$667/A final_adder.U$$666/A VGND VGND VPWR VPWR
+ final_adder.U$$278/B sky130_fd_sc_hd__and2_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3839 _673_/Q U$$3839/B VGND VGND VPWR VPWR U$$3839/X sky130_fd_sc_hd__and2_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_3 dadda_fa_3_31_3/A dadda_fa_3_31_3/B dadda_fa_3_31_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/B dadda_fa_4_31_2/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$183 final_adder.U$$677/A final_adder.U$$549/B1 final_adder.U$$183/B1
+ VGND VGND VPWR VPWR final_adder.U$$183/X sky130_fd_sc_hd__a21o_1
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$194 final_adder.U$$689/A final_adder.U$$688/A VGND VGND VPWR VPWR
+ final_adder.U$$288/A sky130_fd_sc_hd__and2_1
XFILLER_166_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ _543_/CLK _524_/D VGND VGND VPWR VPWR _524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_24_2 U$$1518/X U$$1651/X U$$1727/B VGND VGND VPWR VPWR dadda_fa_4_25_1/A
+ dadda_fa_4_24_2/B sky130_fd_sc_hd__fa_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _455_/CLK _455_/D VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_386_ _515_/CLK _386_/D VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_76_5 dadda_fa_2_76_5/A dadda_fa_2_76_5/B dadda_fa_2_76_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_2/A dadda_fa_4_76_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_69_4 dadda_fa_2_69_4/A dadda_fa_2_69_4/B dadda_fa_2_69_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/CIN dadda_fa_3_69_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_1_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 c[3] VGND VGND VPWR VPWR input190/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_724__776 VGND VGND VPWR VPWR _724__776/HI U$$1787/A1 sky130_fd_sc_hd__conb_1
XFILLER_17_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_106_1 dadda_fa_5_106_1/A dadda_fa_5_106_1/B dadda_fa_5_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/B dadda_fa_7_106_0/A sky130_fd_sc_hd__fa_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_71_4 U$$3740/X U$$3873/X U$$4006/X VGND VGND VPWR VPWR dadda_fa_2_72_1/CIN
+ dadda_fa_2_71_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_64_3 U$$3726/X U$$3859/X U$$3992/X VGND VGND VPWR VPWR dadda_fa_2_65_1/B
+ dadda_fa_2_64_4/B sky130_fd_sc_hd__fa_1
XFILLER_28_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_41_2 dadda_fa_4_41_2/A dadda_fa_4_41_2/B dadda_fa_4_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/CIN dadda_fa_5_41_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_57_2 U$$1983/X U$$2116/X U$$2249/X VGND VGND VPWR VPWR dadda_fa_2_58_1/A
+ dadda_fa_2_57_4/A sky130_fd_sc_hd__fa_1
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_34_1 dadda_fa_4_34_1/A dadda_fa_4_34_1/B dadda_fa_4_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/B dadda_fa_5_34_1/B sky130_fd_sc_hd__fa_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_11_0 dadda_fa_7_11_0/A dadda_fa_7_11_0/B dadda_fa_7_11_0/CIN VGND VGND
+ VPWR VPWR _436_/D _307_/D sky130_fd_sc_hd__fa_2
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_27_0 dadda_fa_4_27_0/A dadda_fa_4_27_0/B dadda_fa_4_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/A dadda_fa_5_27_1/A sky130_fd_sc_hd__fa_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_240_ _499_/CLK _240_/D VGND VGND VPWR VPWR _240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_171_ _448_/CLK _171_/D VGND VGND VPWR VPWR _171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_60_4 U$$1723/X U$$1856/X VGND VGND VPWR VPWR dadda_fa_1_61_7/B dadda_fa_2_60_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_112_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_79_3 dadda_fa_3_79_3/A dadda_fa_3_79_3/B dadda_fa_3_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/B dadda_fa_4_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4304 U$$4304/A U$$4332/B VGND VGND VPWR VPWR U$$4304/X sky130_fd_sc_hd__xor2_1
XU$$4315 _582_/Q U$$4377/A2 U$$70/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4316/A sky130_fd_sc_hd__a22o_1
XU$$4326 U$$4326/A U$$4332/B VGND VGND VPWR VPWR U$$4326/X sky130_fd_sc_hd__xor2_1
XU$$4337 U$$90/A1 U$$4381/A2 U$$4476/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4338/A sky130_fd_sc_hd__a22o_1
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
XU$$4348 U$$4348/A U$$4384/A VGND VGND VPWR VPWR U$$4348/X sky130_fd_sc_hd__xor2_1
XFILLER_93_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3603 U$$3603/A U$$3625/B VGND VGND VPWR VPWR U$$3603/X sky130_fd_sc_hd__xor2_1
XU$$4359 U$$4496/A1 U$$4377/A2 _605_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4360/A sky130_fd_sc_hd__a22o_1
XU$$3614 _574_/Q U$$3678/A2 U$$4438/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3615/A sky130_fd_sc_hd__a22o_1
XFILLER_46_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3625 U$$3625/A U$$3625/B VGND VGND VPWR VPWR U$$3625/X sky130_fd_sc_hd__xor2_1
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3636 U$$4045/B1 U$$3678/A2 U$$76/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3637/A sky130_fd_sc_hd__a22o_1
XU$$2902 U$$2902/A U$$2996/B VGND VGND VPWR VPWR U$$2902/X sky130_fd_sc_hd__xor2_1
XU$$3647 U$$3647/A U$$3699/A VGND VGND VPWR VPWR U$$3647/X sky130_fd_sc_hd__xor2_1
XFILLER_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2913 U$$4283/A1 U$$2975/A2 U$$4285/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2914/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3658 _596_/Q U$$3668/A2 _597_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3659/A sky130_fd_sc_hd__a22o_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2924 U$$2924/A U$$2996/B VGND VGND VPWR VPWR U$$2924/X sky130_fd_sc_hd__xor2_1
XU$$3669 U$$3669/A U$$3699/A VGND VGND VPWR VPWR U$$3669/X sky130_fd_sc_hd__xor2_1
XU$$2935 U$$880/A1 U$$2975/A2 _578_/Q U$$2975/B2 VGND VGND VPWR VPWR U$$2936/A sky130_fd_sc_hd__a22o_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2946 U$$2946/A U$$3004/B VGND VGND VPWR VPWR U$$2946/X sky130_fd_sc_hd__xor2_1
XFILLER_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2957 U$$80/A1 U$$2975/A2 U$$630/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2958/A sky130_fd_sc_hd__a22o_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2968 U$$2968/A U$$3004/B VGND VGND VPWR VPWR U$$2968/X sky130_fd_sc_hd__xor2_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ _510_/CLK _507_/D VGND VGND VPWR VPWR _507_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2979 U$$924/A1 U$$2881/X _600_/Q U$$2882/X VGND VGND VPWR VPWR U$$2980/A sky130_fd_sc_hd__a22o_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _438_/CLK _438_/D VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_369_ _369_/CLK _369_/D VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_81_3 dadda_fa_2_81_3/A dadda_fa_2_81_3/B dadda_fa_2_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/B dadda_fa_3_81_3/B sky130_fd_sc_hd__fa_1
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_2 dadda_fa_2_74_2/A dadda_fa_2_74_2/B dadda_fa_2_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/A dadda_fa_3_74_3/A sky130_fd_sc_hd__fa_2
XFILLER_111_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_51_1 dadda_fa_5_51_1/A dadda_fa_5_51_1/B dadda_fa_5_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/B dadda_fa_7_51_0/A sky130_fd_sc_hd__fa_1
XFILLER_123_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_67_1 dadda_fa_2_67_1/A dadda_fa_2_67_1/B dadda_fa_2_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/CIN dadda_fa_3_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_44_0 dadda_fa_5_44_0/A dadda_fa_5_44_0/B dadda_fa_5_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/A dadda_fa_6_44_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_96_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_89_2 dadda_fa_4_89_2/A dadda_fa_4_89_2/B dadda_fa_4_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/CIN dadda_fa_5_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_59_0 dadda_fa_7_59_0/A dadda_fa_7_59_0/B dadda_fa_7_59_0/CIN VGND VGND
+ VPWR VPWR _484_/D _355_/D sky130_fd_sc_hd__fa_2
XFILLER_154_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_62_0 U$$2392/X U$$2525/X U$$2658/X VGND VGND VPWR VPWR dadda_fa_2_63_0/B
+ dadda_fa_2_62_3/B sky130_fd_sc_hd__fa_2
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2209 U$$2209/A U$$2289/B VGND VGND VPWR VPWR U$$2209/X sky130_fd_sc_hd__xor2_1
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1508 _638_/Q VGND VGND VPWR VPWR U$$1510/B sky130_fd_sc_hd__inv_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1519 U$$971/A1 U$$1511/X U$$12/B1 U$$1512/X VGND VGND VPWR VPWR U$$1520/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_223_ _474_/CLK _223_/D VGND VGND VPWR VPWR _223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_91_2 dadda_fa_3_91_2/A dadda_fa_3_91_2/B dadda_fa_3_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/A dadda_fa_4_91_2/B sky130_fd_sc_hd__fa_2
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_84_1 dadda_fa_3_84_1/A dadda_fa_3_84_1/B dadda_fa_3_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/CIN dadda_fa_4_84_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_61_0 dadda_fa_6_61_0/A dadda_fa_6_61_0/B dadda_fa_6_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_62_0/B dadda_fa_7_61_0/CIN sky130_fd_sc_hd__fa_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_77_0 dadda_fa_3_77_0/A dadda_fa_3_77_0/B dadda_fa_3_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/B dadda_fa_4_77_1/CIN sky130_fd_sc_hd__fa_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater408 U$$3545/A2 VGND VGND VPWR VPWR U$$3525/A2 sky130_fd_sc_hd__buf_12
XFILLER_120_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4101 U$$539/A1 U$$4107/A2 _613_/Q U$$4107/B2 VGND VGND VPWR VPWR U$$4102/A sky130_fd_sc_hd__a22o_1
Xrepeater419 U$$2870/A2 VGND VGND VPWR VPWR U$$2868/A2 sky130_fd_sc_hd__buf_12
XU$$4112 U$$4197/B VGND VGND VPWR VPWR U$$4112/Y sky130_fd_sc_hd__inv_1
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4123 U$$4123/A U$$4197/B VGND VGND VPWR VPWR U$$4123/X sky130_fd_sc_hd__xor2_1
XFILLER_66_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4134 U$$4271/A1 U$$4114/X U$$4273/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4135/A
+ sky130_fd_sc_hd__a22o_1
XU$$4145 U$$4145/A _677_/Q VGND VGND VPWR VPWR U$$4145/X sky130_fd_sc_hd__xor2_1
XU$$3400 U$$4496/A1 U$$3292/X _605_/Q U$$3293/X VGND VGND VPWR VPWR U$$3401/A sky130_fd_sc_hd__a22o_1
XFILLER_93_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3411 U$$3411/A U$$3413/B VGND VGND VPWR VPWR U$$3411/X sky130_fd_sc_hd__xor2_1
XU$$4156 U$$4291/B1 U$$4114/X U$$4156/B1 U$$4198/B2 VGND VGND VPWR VPWR U$$4157/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_113_1 input144/X dadda_fa_4_113_1/B dadda_fa_4_113_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_114_0/B dadda_fa_5_113_1/B sky130_fd_sc_hd__fa_1
XU$$3422 U$$819/A1 U$$3292/X U$$3422/B1 U$$3293/X VGND VGND VPWR VPWR U$$3423/A sky130_fd_sc_hd__a22o_1
XU$$4167 U$$4167/A U$$4247/A VGND VGND VPWR VPWR U$$4167/X sky130_fd_sc_hd__xor2_1
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4178 U$$4178/A1 U$$4114/X U$$70/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4179/A sky130_fd_sc_hd__a22o_1
XU$$3433 U$$4255/A1 U$$3525/A2 _553_/Q U$$3525/B2 VGND VGND VPWR VPWR U$$3434/A sky130_fd_sc_hd__a22o_1
XU$$3444 U$$3444/A U$$3561/A VGND VGND VPWR VPWR U$$3444/X sky130_fd_sc_hd__xor2_1
XU$$4189 U$$4189/A U$$4247/A VGND VGND VPWR VPWR U$$4189/X sky130_fd_sc_hd__xor2_1
XU$$2710 U$$2710/A U$$2710/B VGND VGND VPWR VPWR U$$2710/X sky130_fd_sc_hd__xor2_1
XU$$3455 U$$30/A1 U$$3525/A2 U$$30/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3456/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_0 dadda_fa_4_106_0/A dadda_fa_4_106_0/B dadda_fa_4_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/A dadda_fa_5_106_1/A sky130_fd_sc_hd__fa_1
XU$$2721 U$$940/A1 U$$2729/A2 U$$942/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2722/A sky130_fd_sc_hd__a22o_1
XU$$3466 U$$3466/A _667_/Q VGND VGND VPWR VPWR U$$3466/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_39_5 dadda_fa_2_39_5/A dadda_fa_2_39_5/B dadda_fa_2_39_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_40_2/A dadda_fa_4_39_0/A sky130_fd_sc_hd__fa_1
XFILLER_19_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2732 U$$2732/A _655_/Q VGND VGND VPWR VPWR U$$2732/X sky130_fd_sc_hd__xor2_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3477 _574_/Q U$$3545/A2 _575_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3478/A sky130_fd_sc_hd__a22o_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3488 U$$3488/A U$$3496/B VGND VGND VPWR VPWR U$$3488/X sky130_fd_sc_hd__xor2_1
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2743 _657_/Q U$$2743/B VGND VGND VPWR VPWR U$$2743/X sky130_fd_sc_hd__and2_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3499 _585_/Q U$$3545/A2 _586_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3500/A sky130_fd_sc_hd__a22o_1
XU$$2754 U$$14/A1 U$$2796/A2 _556_/Q U$$2826/B2 VGND VGND VPWR VPWR U$$2755/A sky130_fd_sc_hd__a22o_1
XU$$2765 U$$2765/A U$$2797/B VGND VGND VPWR VPWR U$$2765/X sky130_fd_sc_hd__xor2_1
XU$$2776 U$$36/A1 U$$2796/A2 _567_/Q U$$2745/X VGND VGND VPWR VPWR U$$2777/A sky130_fd_sc_hd__a22o_1
XU$$2787 U$$2787/A U$$2839/B VGND VGND VPWR VPWR U$$2787/X sky130_fd_sc_hd__xor2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2798 U$$58/A1 U$$2868/A2 _578_/Q U$$2745/X VGND VGND VPWR VPWR U$$2799/A sky130_fd_sc_hd__a22o_1
X_795__847 VGND VGND VPWR VPWR _795__847/HI U$$4435/B sky130_fd_sc_hd__conb_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_836__888 VGND VGND VPWR VPWR _836__888/HI U$$4517/B sky130_fd_sc_hd__conb_1
Xdadda_fa_5_99_1 dadda_fa_5_99_1/A dadda_fa_5_99_1/B dadda_fa_5_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/B dadda_fa_7_99_0/A sky130_fd_sc_hd__fa_2
XFILLER_105_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$705 final_adder.U$$705/A final_adder.U$$705/B VGND VGND VPWR VPWR
+ _251_/D sky130_fd_sc_hd__xor2_1
XFILLER_151_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$716 final_adder.U$$716/A final_adder.U$$716/B VGND VGND VPWR VPWR
+ _262_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$727 final_adder.U$$727/A final_adder.U$$727/B VGND VGND VPWR VPWR
+ _273_/D sky130_fd_sc_hd__xor2_1
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$738 final_adder.U$$738/A final_adder.U$$738/B VGND VGND VPWR VPWR
+ _284_/D sky130_fd_sc_hd__xor2_1
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$749 final_adder.U$$749/A final_adder.U$$749/B VGND VGND VPWR VPWR
+ _295_/D sky130_fd_sc_hd__xor2_2
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_94_0 dadda_fa_4_94_0/A dadda_fa_4_94_0/B dadda_fa_4_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/A dadda_fa_5_94_1/A sky130_fd_sc_hd__fa_1
XFILLER_193_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_108_2 U$$4080/X U$$4213/X U$$4346/X VGND VGND VPWR VPWR dadda_fa_4_109_1/A
+ dadda_fa_4_108_2/B sky130_fd_sc_hd__fa_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput280 _288_/Q VGND VGND VPWR VPWR o[120] sky130_fd_sc_hd__buf_2
Xoutput291 _183_/Q VGND VGND VPWR VPWR o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2006 U$$771/B1 U$$2052/A2 U$$912/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2007/A sky130_fd_sc_hd__a22o_1
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2017 U$$2017/A U$$2023/B VGND VGND VPWR VPWR U$$2017/X sky130_fd_sc_hd__xor2_1
XFILLER_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2028 U$$932/A1 U$$2052/A2 U$$934/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2029/A sky130_fd_sc_hd__a22o_1
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2039 U$$2039/A U$$2055/A VGND VGND VPWR VPWR U$$2039/X sky130_fd_sc_hd__xor2_1
XFILLER_43_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1305 U$$892/B1 U$$1367/A2 U$$74/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1306/A sky130_fd_sc_hd__a22o_1
XU$$1316 U$$1316/A U$$1369/A VGND VGND VPWR VPWR U$$1316/X sky130_fd_sc_hd__xor2_1
XU$$1327 U$$92/B1 U$$1341/A2 U$$96/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1328/A sky130_fd_sc_hd__a22o_1
XU$$1338 U$$1338/A U$$1369/A VGND VGND VPWR VPWR U$$1338/X sky130_fd_sc_hd__xor2_1
XU$$1349 U$$938/A1 U$$1367/A2 U$$940/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1350/A sky130_fd_sc_hd__a22o_1
XFILLER_70_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ _448_/CLK _206_/D VGND VGND VPWR VPWR _206_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_51_4 dadda_fa_2_51_4/A dadda_fa_2_51_4/B dadda_fa_2_51_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/CIN dadda_fa_3_51_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_44_3 dadda_fa_2_44_3/A dadda_fa_2_44_3/B dadda_fa_2_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/B dadda_fa_3_44_3/B sky130_fd_sc_hd__fa_1
XU$$3230 U$$3230/A U$$3244/B VGND VGND VPWR VPWR U$$3230/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$12 _436_/Q _308_/Q VGND VGND VPWR VPWR final_adder.U$$507/B1 final_adder.U$$634/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3241 U$$912/A1 U$$3241/A2 U$$4476/A1 U$$3253/B2 VGND VGND VPWR VPWR U$$3242/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$23 _447_/Q _319_/Q VGND VGND VPWR VPWR final_adder.U$$151/B1 final_adder.U$$645/A
+ sky130_fd_sc_hd__ha_1
XFILLER_111_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$34 _458_/Q _330_/Q VGND VGND VPWR VPWR final_adder.U$$529/B1 final_adder.U$$656/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_2 U$$1544/X U$$1677/X U$$1810/X VGND VGND VPWR VPWR dadda_fa_3_38_1/A
+ dadda_fa_3_37_3/A sky130_fd_sc_hd__fa_1
XU$$3252 U$$3252/A _663_/Q VGND VGND VPWR VPWR U$$3252/X sky130_fd_sc_hd__xor2_1
XU$$3263 U$$4496/A1 U$$3155/X _605_/Q U$$3156/X VGND VGND VPWR VPWR U$$3264/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$45 _469_/Q _341_/Q VGND VGND VPWR VPWR final_adder.U$$173/B1 final_adder.U$$667/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3274 U$$3274/A _663_/Q VGND VGND VPWR VPWR U$$3274/X sky130_fd_sc_hd__xor2_1
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$56 _480_/Q _352_/Q VGND VGND VPWR VPWR final_adder.U$$551/B1 final_adder.U$$678/A
+ sky130_fd_sc_hd__ha_1
XU$$2540 U$$4045/B1 U$$2584/A2 _586_/Q U$$2584/B2 VGND VGND VPWR VPWR U$$2541/A sky130_fd_sc_hd__a22o_1
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3285 U$$956/A1 U$$3155/X U$$3285/B1 U$$3156/X VGND VGND VPWR VPWR U$$3286/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$67 _491_/Q _363_/Q VGND VGND VPWR VPWR final_adder.U$$195/B1 final_adder.U$$689/A
+ sky130_fd_sc_hd__ha_1
XU$$2551 U$$2551/A U$$2585/B VGND VGND VPWR VPWR U$$2551/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_1 dadda_fa_5_14_1/A dadda_fa_5_14_1/B dadda_fa_5_14_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/B dadda_fa_7_14_0/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$78 _502_/Q _374_/Q VGND VGND VPWR VPWR final_adder.U$$573/B1 final_adder.U$$700/A
+ sky130_fd_sc_hd__ha_1
XFILLER_59_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3296 U$$4255/A1 U$$3412/A2 U$$969/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3297/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2562 U$$96/A1 U$$2584/A2 U$$96/B1 U$$2584/B2 VGND VGND VPWR VPWR U$$2563/A sky130_fd_sc_hd__a22o_1
XFILLER_179_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$89 _513_/Q _385_/Q VGND VGND VPWR VPWR final_adder.U$$217/B1 final_adder.U$$711/A
+ sky130_fd_sc_hd__ha_1
XU$$2573 U$$2573/A U$$2603/A VGND VGND VPWR VPWR U$$2573/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2584 _607_/Q U$$2584/A2 _608_/Q U$$2584/B2 VGND VGND VPWR VPWR U$$2585/A sky130_fd_sc_hd__a22o_1
XFILLER_181_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1850 U$$1850/A U$$1856/B VGND VGND VPWR VPWR U$$1850/X sky130_fd_sc_hd__xor2_1
XU$$2595 U$$2595/A _653_/Q VGND VGND VPWR VPWR U$$2595/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1861 U$$80/A1 U$$1785/X U$$82/A1 U$$1786/X VGND VGND VPWR VPWR U$$1862/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1872 U$$1872/A U$$1872/B VGND VGND VPWR VPWR U$$1872/X sky130_fd_sc_hd__xor2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1883 _599_/Q U$$1903/A2 _600_/Q U$$1903/B2 VGND VGND VPWR VPWR U$$1884/A sky130_fd_sc_hd__a22o_1
XU$$1894 U$$1894/A _643_/Q VGND VGND VPWR VPWR U$$1894/X sky130_fd_sc_hd__xor2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$513 final_adder.U$$640/A final_adder.U$$640/B final_adder.U$$513/B1
+ VGND VGND VPWR VPWR final_adder.U$$641/B sky130_fd_sc_hd__a21o_1
XFILLER_9_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$535 final_adder.U$$662/A final_adder.U$$662/B final_adder.U$$535/B1
+ VGND VGND VPWR VPWR final_adder.U$$663/B sky130_fd_sc_hd__a21o_1
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater750 _557_/Q VGND VGND VPWR VPWR U$$4265/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$557 final_adder.U$$684/A final_adder.U$$684/B final_adder.U$$557/B1
+ VGND VGND VPWR VPWR final_adder.U$$685/B sky130_fd_sc_hd__a21o_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater761 _552_/Q VGND VGND VPWR VPWR U$$4255/A1 sky130_fd_sc_hd__buf_12
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$407 U$$407/A _621_/Q VGND VGND VPWR VPWR U$$407/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$579 final_adder.U$$706/A final_adder.U$$706/B final_adder.U$$579/B1
+ VGND VGND VPWR VPWR final_adder.U$$707/B sky130_fd_sc_hd__a21o_1
XU$$418 U$$418/A U$$547/A VGND VGND VPWR VPWR U$$418/X sky130_fd_sc_hd__xor2_1
XU$$429 U$$18/A1 U$$491/A2 U$$20/A1 U$$416/X VGND VGND VPWR VPWR U$$430/A sky130_fd_sc_hd__a22o_1
XFILLER_44_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_113_0 U$$3424/Y U$$3558/X U$$3691/X VGND VGND VPWR VPWR dadda_fa_4_114_1/CIN
+ dadda_fa_4_113_2/B sky130_fd_sc_hd__fa_1
XFILLER_119_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_61_3 dadda_fa_3_61_3/A dadda_fa_3_61_3/B dadda_fa_3_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/B dadda_fa_4_61_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_54_2 dadda_fa_3_54_2/A dadda_fa_3_54_2/B dadda_fa_3_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/A dadda_fa_4_54_2/B sky130_fd_sc_hd__fa_2
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_47_1 dadda_fa_3_47_1/A dadda_fa_3_47_1/B dadda_fa_3_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/CIN dadda_fa_4_47_2/A sky130_fd_sc_hd__fa_1
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_24_0 dadda_fa_6_24_0/A dadda_fa_6_24_0/B dadda_fa_6_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_25_0/B dadda_fa_7_24_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$930 U$$930/A1 U$$826/X U$$932/A1 U$$827/X VGND VGND VPWR VPWR U$$931/A sky130_fd_sc_hd__a22o_1
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$941 U$$941/A U$$943/B VGND VGND VPWR VPWR U$$941/X sky130_fd_sc_hd__xor2_1
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$952 U$$952/A1 U$$826/X U$$952/B1 U$$827/X VGND VGND VPWR VPWR U$$953/A sky130_fd_sc_hd__a22o_1
XFILLER_44_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1102 U$$1102/A1 U$$1100/X _552_/Q U$$1101/X VGND VGND VPWR VPWR U$$1103/A sky130_fd_sc_hd__a22o_1
XU$$963 U$$961/Y _630_/Q U$$959/A U$$962/X U$$959/Y VGND VGND VPWR VPWR U$$963/X sky130_fd_sc_hd__a32o_4
XFILLER_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$974 U$$974/A U$$992/B VGND VGND VPWR VPWR U$$974/X sky130_fd_sc_hd__xor2_1
XU$$1113 U$$1113/A U$$1167/B VGND VGND VPWR VPWR U$$1113/X sky130_fd_sc_hd__xor2_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1124 U$$987/A1 U$$1200/A2 U$$28/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1125/A sky130_fd_sc_hd__a22o_1
XU$$985 U$$26/A1 U$$999/A2 U$$987/A1 U$$987/B2 VGND VGND VPWR VPWR U$$986/A sky130_fd_sc_hd__a22o_1
XU$$996 U$$996/A U$$998/B VGND VGND VPWR VPWR U$$996/X sky130_fd_sc_hd__xor2_1
XU$$1135 U$$1135/A U$$1167/B VGND VGND VPWR VPWR U$$1135/X sky130_fd_sc_hd__xor2_1
XU$$1146 U$$50/A1 U$$1200/A2 U$$50/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1147/A sky130_fd_sc_hd__a22o_1
XFILLER_71_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1157 U$$1157/A U$$1167/B VGND VGND VPWR VPWR U$$1157/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_112_2 U$$4088/X U$$4221/X VGND VGND VPWR VPWR dadda_fa_4_113_2/A dadda_ha_3_112_2/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1168 U$$72/A1 U$$1218/A2 U$$74/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1169/A sky130_fd_sc_hd__a22o_1
XU$$1179 U$$1179/A U$$1232/A VGND VGND VPWR VPWR U$$1179/X sky130_fd_sc_hd__xor2_1
XFILLER_31_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_99_4 U$$4062/X U$$4195/X U$$4328/X VGND VGND VPWR VPWR dadda_fa_3_100_2/B
+ dadda_fa_4_99_0/A sky130_fd_sc_hd__fa_1
XFILLER_172_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_42_0 U$$1953/X U$$2086/X U$$2219/X VGND VGND VPWR VPWR dadda_fa_3_43_0/B
+ dadda_fa_3_42_2/B sky130_fd_sc_hd__fa_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3060 U$$46/A1 U$$3146/A2 _572_/Q U$$3146/B2 VGND VGND VPWR VPWR U$$3061/A sky130_fd_sc_hd__a22o_1
XU$$3071 U$$3071/A U$$3085/B VGND VGND VPWR VPWR U$$3071/X sky130_fd_sc_hd__xor2_1
XFILLER_179_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3082 U$$4178/A1 U$$3146/A2 U$$892/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3083/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3093 U$$3093/A U$$3109/B VGND VGND VPWR VPWR U$$3093/X sky130_fd_sc_hd__xor2_1
XU$$2370 U$$2370/A U$$2436/B VGND VGND VPWR VPWR U$$2370/X sky130_fd_sc_hd__xor2_1
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2381 U$$50/B1 U$$2421/A2 U$$4438/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2382/A sky130_fd_sc_hd__a22o_1
XFILLER_50_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2392 U$$2392/A U$$2432/B VGND VGND VPWR VPWR U$$2392/X sky130_fd_sc_hd__xor2_1
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1680 U$$36/A1 U$$1734/A2 U$$38/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1681/A sky130_fd_sc_hd__a22o_1
XU$$1691 U$$1691/A U$$1739/B VGND VGND VPWR VPWR U$$1691/X sky130_fd_sc_hd__xor2_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_88_4 U$$3242/X U$$3375/X VGND VGND VPWR VPWR dadda_fa_2_89_4/CIN dadda_fa_3_88_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_120_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_71_2 dadda_fa_4_71_2/A dadda_fa_4_71_2/B dadda_fa_4_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/CIN dadda_fa_5_71_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_2 U$$2442/X U$$2575/X U$$2708/X VGND VGND VPWR VPWR dadda_fa_2_88_3/CIN
+ dadda_fa_2_87_5/B sky130_fd_sc_hd__fa_1
XFILLER_143_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_64_1 dadda_fa_4_64_1/A dadda_fa_4_64_1/B dadda_fa_4_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/B dadda_fa_5_64_1/B sky130_fd_sc_hd__fa_1
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_41_0 dadda_fa_7_41_0/A dadda_fa_7_41_0/B dadda_fa_7_41_0/CIN VGND VGND
+ VPWR VPWR _466_/D _337_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_57_0 dadda_fa_4_57_0/A dadda_fa_4_57_0/B dadda_fa_4_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/A dadda_fa_5_57_1/A sky130_fd_sc_hd__fa_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$310 final_adder.U$$310/A final_adder.U$$310/B VGND VGND VPWR VPWR
+ final_adder.U$$346/A sky130_fd_sc_hd__and2_1
XFILLER_188_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$321 final_adder.U$$258/X final_adder.U$$626/B final_adder.U$$259/X
+ VGND VGND VPWR VPWR final_adder.U$$630/B sky130_fd_sc_hd__a21o_2
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$332 final_adder.U$$332/A final_adder.U$$332/B VGND VGND VPWR VPWR
+ final_adder.U$$358/B sky130_fd_sc_hd__and2_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$343 final_adder.U$$342/A final_adder.U$$301/X final_adder.U$$303/X
+ VGND VGND VPWR VPWR final_adder.U$$343/X sky130_fd_sc_hd__a21o_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$354 final_adder.U$$354/A final_adder.U$$354/B VGND VGND VPWR VPWR
+ final_adder.U$$354/X sky130_fd_sc_hd__and2_1
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$365 final_adder.U$$364/A final_adder.U$$345/X final_adder.U$$347/X
+ VGND VGND VPWR VPWR final_adder.U$$365/X sky130_fd_sc_hd__a21o_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$204 U$$204/A U$$274/A VGND VGND VPWR VPWR U$$204/X sky130_fd_sc_hd__xor2_1
XFILLER_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$215 U$$78/A1 U$$141/X U$$80/A1 U$$142/X VGND VGND VPWR VPWR U$$216/A sky130_fd_sc_hd__a22o_1
Xrepeater580 _639_/Q VGND VGND VPWR VPWR U$$1643/A sky130_fd_sc_hd__buf_12
XFILLER_85_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_540_ _543_/CLK _540_/D VGND VGND VPWR VPWR _540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$387 final_adder.U$$372/B final_adder.U$$686/B final_adder.U$$361/X
+ VGND VGND VPWR VPWR final_adder.U$$702/B sky130_fd_sc_hd__a21o_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$226 U$$226/A U$$242/B VGND VGND VPWR VPWR U$$226/X sky130_fd_sc_hd__xor2_1
Xrepeater591 _631_/Q VGND VGND VPWR VPWR U$$980/B sky130_fd_sc_hd__buf_12
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$237 U$$98/B1 U$$141/X U$$924/A1 U$$142/X VGND VGND VPWR VPWR U$$238/A sky130_fd_sc_hd__a22o_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$248 U$$248/A U$$262/B VGND VGND VPWR VPWR U$$248/X sky130_fd_sc_hd__xor2_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$259 U$$944/A1 U$$141/X U$$946/A1 U$$142/X VGND VGND VPWR VPWR U$$260/A sky130_fd_sc_hd__a22o_1
XFILLER_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ _471_/CLK _471_/D VGND VGND VPWR VPWR _471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$9 U$$9/A U$$9/B VGND VGND VPWR VPWR U$$9/X sky130_fd_sc_hd__xor2_2
XFILLER_5_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_75_0 U$$821/Y U$$955/X U$$1088/X VGND VGND VPWR VPWR dadda_fa_1_76_8/A
+ dadda_fa_1_75_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$760 U$$760/A U$$784/B VGND VGND VPWR VPWR U$$760/X sky130_fd_sc_hd__xor2_1
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_669_ _669_/CLK _669_/D VGND VGND VPWR VPWR _669_/Q sky130_fd_sc_hd__dfxtp_4
XU$$771 U$$771/A1 U$$689/X U$$771/B1 U$$690/X VGND VGND VPWR VPWR U$$772/A sky130_fd_sc_hd__a22o_1
XU$$782 U$$782/A _627_/Q VGND VGND VPWR VPWR U$$782/X sky130_fd_sc_hd__xor2_2
XU$$793 U$$928/B1 U$$817/A2 _603_/Q U$$817/B2 VGND VGND VPWR VPWR U$$794/A sky130_fd_sc_hd__a22o_1
XFILLER_189_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_81_1 dadda_fa_5_81_1/A dadda_fa_5_81_1/B dadda_fa_5_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/B dadda_fa_7_81_0/A sky130_fd_sc_hd__fa_1
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_97_1 U$$2728/X U$$2861/X U$$2994/X VGND VGND VPWR VPWR dadda_fa_3_98_0/CIN
+ dadda_fa_3_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_74_0 dadda_fa_5_74_0/A dadda_fa_5_74_0/B dadda_fa_5_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/A dadda_fa_6_74_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_73_8 dadda_fa_1_73_8/A dadda_fa_1_73_8/B dadda_fa_1_73_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_3/A dadda_fa_3_73_0/A sky130_fd_sc_hd__fa_2
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_66_7 dadda_fa_1_66_7/A dadda_fa_1_66_7/B dadda_fa_1_66_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/CIN dadda_fa_2_66_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_6 U$$3982/X input211/X dadda_fa_1_59_6/CIN VGND VGND VPWR VPWR dadda_fa_2_60_2/B
+ dadda_fa_2_59_5/B sky130_fd_sc_hd__fa_2
XFILLER_187_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_89_0 dadda_fa_7_89_0/A dadda_fa_7_89_0/B dadda_fa_7_89_0/CIN VGND VGND
+ VPWR VPWR _514_/D _385_/D sky130_fd_sc_hd__fa_2
XFILLER_175_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_92_0 _691__911/HI U$$2053/X U$$2186/X VGND VGND VPWR VPWR dadda_fa_2_93_4/CIN
+ dadda_fa_2_92_5/B sky130_fd_sc_hd__fa_2
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4508 U$$4508/A1 U$$4388/X U$$4510/A1 U$$4389/X VGND VGND VPWR VPWR U$$4509/A sky130_fd_sc_hd__a22o_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$140 final_adder.U$$635/A final_adder.U$$634/A VGND VGND VPWR VPWR
+ final_adder.U$$262/B sky130_fd_sc_hd__and2_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3807 U$$4492/A1 U$$3703/X U$$4494/A1 U$$3704/X VGND VGND VPWR VPWR U$$3808/A sky130_fd_sc_hd__a22o_1
XFILLER_131_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3818 U$$3818/A U$$3835/A VGND VGND VPWR VPWR U$$3818/X sky130_fd_sc_hd__xor2_1
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$151 final_adder.U$$645/A final_adder.U$$517/B1 final_adder.U$$151/B1
+ VGND VGND VPWR VPWR final_adder.U$$151/X sky130_fd_sc_hd__a21o_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3829 _613_/Q U$$3703/X U$$4379/A1 U$$3704/X VGND VGND VPWR VPWR U$$3830/A sky130_fd_sc_hd__a22o_1
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$162 final_adder.U$$657/A final_adder.U$$656/A VGND VGND VPWR VPWR
+ final_adder.U$$272/A sky130_fd_sc_hd__and2_1
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_104_0 dadda_fa_6_104_0/A dadda_fa_6_104_0/B dadda_fa_6_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_105_0/B dadda_fa_7_104_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$173 final_adder.U$$667/A final_adder.U$$539/B1 final_adder.U$$173/B1
+ VGND VGND VPWR VPWR final_adder.U$$173/X sky130_fd_sc_hd__a21o_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$184 final_adder.U$$679/A final_adder.U$$678/A VGND VGND VPWR VPWR
+ final_adder.U$$284/B sky130_fd_sc_hd__and2_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$195 final_adder.U$$689/A final_adder.U$$561/B1 final_adder.U$$195/B1
+ VGND VGND VPWR VPWR final_adder.U$$195/X sky130_fd_sc_hd__a21o_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_523_ _583_/CLK _523_/D VGND VGND VPWR VPWR _523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_24_3 input173/X dadda_fa_3_24_3/B dadda_fa_3_24_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_25_1/B dadda_fa_4_24_2/CIN sky130_fd_sc_hd__fa_2
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ _454_/CLK _454_/D VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_385_ _518_/CLK _385_/D VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_91_0 dadda_fa_6_91_0/A dadda_fa_6_91_0/B dadda_fa_6_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_92_0/B dadda_fa_7_91_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_127_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_69_5 dadda_fa_2_69_5/A dadda_fa_2_69_5/B dadda_fa_2_69_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_2/A dadda_fa_4_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_1_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput180 c[30] VGND VGND VPWR VPWR input180/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput191 c[40] VGND VGND VPWR VPWR input191/X sky130_fd_sc_hd__buf_2
XFILLER_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$590 _569_/Q U$$626/A2 _570_/Q U$$553/X VGND VGND VPWR VPWR U$$591/A sky130_fd_sc_hd__a22o_1
XFILLER_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_71_5 U$$4139/X U$$4272/X U$$4405/X VGND VGND VPWR VPWR dadda_fa_2_72_2/A
+ dadda_fa_2_71_5/A sky130_fd_sc_hd__fa_1
XFILLER_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_64_4 U$$4125/X U$$4258/X U$$4391/X VGND VGND VPWR VPWR dadda_fa_2_65_1/CIN
+ dadda_fa_2_64_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_189_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_3 U$$2382/X U$$2515/X U$$2648/X VGND VGND VPWR VPWR dadda_fa_2_58_1/B
+ dadda_fa_2_57_4/B sky130_fd_sc_hd__fa_1
XFILLER_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_34_2 dadda_fa_4_34_2/A dadda_fa_4_34_2/B dadda_fa_4_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/CIN dadda_fa_5_34_1/CIN sky130_fd_sc_hd__fa_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_27_1 dadda_fa_4_27_1/A dadda_fa_4_27_1/B dadda_fa_4_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/B dadda_fa_5_27_1/B sky130_fd_sc_hd__fa_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_170_ _448_/CLK _170_/D VGND VGND VPWR VPWR _170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4305 U$$4442/A1 U$$4377/A2 _578_/Q U$$4377/B2 VGND VGND VPWR VPWR U$$4306/A sky130_fd_sc_hd__a22o_1
XFILLER_120_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4316 U$$4316/A U$$4384/A VGND VGND VPWR VPWR U$$4316/X sky130_fd_sc_hd__xor2_1
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4327 U$$765/A1 U$$4251/X U$$630/A1 U$$4252/X VGND VGND VPWR VPWR U$$4328/A sky130_fd_sc_hd__a22o_1
XU$$4338 U$$4338/A _679_/Q VGND VGND VPWR VPWR U$$4338/X sky130_fd_sc_hd__xor2_1
XU$$3604 U$$4289/A1 U$$3624/A2 U$$4289/B1 U$$3624/B2 VGND VGND VPWR VPWR U$$3605/A
+ sky130_fd_sc_hd__a22o_1
XU$$4349 U$$4486/A1 U$$4381/A2 U$$787/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4350/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_16_1 U$$438/X U$$571/X VGND VGND VPWR VPWR dadda_fa_4_17_2/A dadda_ha_3_16_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3615 U$$3615/A U$$3698/A VGND VGND VPWR VPWR U$$3615/X sky130_fd_sc_hd__xor2_1
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_747__799 VGND VGND VPWR VPWR _747__799/HI U$$3285/B1 sky130_fd_sc_hd__conb_1
XU$$3626 _580_/Q U$$3678/A2 U$$66/A1 U$$3678/B2 VGND VGND VPWR VPWR U$$3627/A sky130_fd_sc_hd__a22o_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3637 U$$3637/A _669_/Q VGND VGND VPWR VPWR U$$3637/X sky130_fd_sc_hd__xor2_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2903 U$$4273/A1 U$$2975/A2 _562_/Q U$$2975/B2 VGND VGND VPWR VPWR U$$2904/A sky130_fd_sc_hd__a22o_1
XU$$3648 _591_/Q U$$3668/A2 U$$4335/A1 U$$3668/B2 VGND VGND VPWR VPWR U$$3649/A sky130_fd_sc_hd__a22o_1
XU$$2914 U$$2914/A U$$2960/B VGND VGND VPWR VPWR U$$2914/X sky130_fd_sc_hd__xor2_1
XU$$3659 U$$3659/A U$$3699/A VGND VGND VPWR VPWR U$$3659/X sky130_fd_sc_hd__xor2_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2925 U$$48/A1 U$$3009/A2 U$$50/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2926/A sky130_fd_sc_hd__a22o_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2936 U$$2936/A U$$2960/B VGND VGND VPWR VPWR U$$2936/X sky130_fd_sc_hd__xor2_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2947 _583_/Q U$$2881/X _584_/Q U$$2882/X VGND VGND VPWR VPWR U$$2948/A sky130_fd_sc_hd__a22o_1
XFILLER_46_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_22_0 U$$317/X U$$450/X U$$583/X VGND VGND VPWR VPWR dadda_fa_4_23_0/B
+ dadda_fa_4_22_1/CIN sky130_fd_sc_hd__fa_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2958 U$$2958/A _659_/Q VGND VGND VPWR VPWR U$$2958/X sky130_fd_sc_hd__xor2_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_506_ _509_/CLK _506_/D VGND VGND VPWR VPWR _506_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2969 U$$4476/A1 U$$2881/X _595_/Q U$$2882/X VGND VGND VPWR VPWR U$$2970/A sky130_fd_sc_hd__a22o_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_437_ _454_/CLK _437_/D VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_368_ _497_/CLK _368_/D VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_299_ _429_/CLK _299_/D VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_81_4 dadda_fa_2_81_4/A dadda_fa_2_81_4/B dadda_fa_2_81_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/CIN dadda_fa_3_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_74_3 dadda_fa_2_74_3/A dadda_fa_2_74_3/B dadda_fa_2_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/B dadda_fa_3_74_3/B sky130_fd_sc_hd__fa_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_67_2 dadda_fa_2_67_2/A dadda_fa_2_67_2/B dadda_fa_2_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/A dadda_fa_3_67_3/A sky130_fd_sc_hd__fa_2
XFILLER_95_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_44_1 dadda_fa_5_44_1/A dadda_fa_5_44_1/B dadda_fa_5_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/B dadda_fa_7_44_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_37_0 dadda_fa_5_37_0/A dadda_fa_5_37_0/B dadda_fa_5_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/A dadda_fa_6_37_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_696__916 VGND VGND VPWR VPWR _696__916/HI _696__916/LO sky130_fd_sc_hd__conb_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_111_0 dadda_fa_5_111_0/A dadda_fa_5_111_0/B dadda_fa_5_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/A dadda_fa_6_111_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_193_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_1 U$$2791/X U$$2924/X U$$3057/X VGND VGND VPWR VPWR dadda_fa_2_63_0/CIN
+ dadda_fa_2_62_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_55_0 U$$782/X U$$915/X U$$1048/X VGND VGND VPWR VPWR dadda_fa_2_56_0/B
+ dadda_fa_2_55_3/B sky130_fd_sc_hd__fa_1
XFILLER_170_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1509 _639_/Q VGND VGND VPWR VPWR U$$1509/Y sky130_fd_sc_hd__inv_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_222_ _480_/CLK _222_/D VGND VGND VPWR VPWR _222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_91_3 dadda_fa_3_91_3/A dadda_fa_3_91_3/B dadda_fa_3_91_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/B dadda_fa_4_91_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_152_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_84_2 dadda_fa_3_84_2/A dadda_fa_3_84_2/B dadda_fa_3_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/A dadda_fa_4_84_2/B sky130_fd_sc_hd__fa_1
XFILLER_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_1 dadda_fa_3_77_1/A dadda_fa_3_77_1/B dadda_fa_3_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/CIN dadda_fa_4_77_2/A sky130_fd_sc_hd__fa_2
XFILLER_152_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_54_0 dadda_fa_6_54_0/A dadda_fa_6_54_0/B dadda_fa_6_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_55_0/B dadda_fa_7_54_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_105_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater409 U$$3429/X VGND VGND VPWR VPWR U$$3545/A2 sky130_fd_sc_hd__buf_12
XU$$4102 U$$4102/A U$$4109/A VGND VGND VPWR VPWR U$$4102/X sky130_fd_sc_hd__xor2_1
XU$$4113 U$$4197/B U$$4113/B VGND VGND VPWR VPWR U$$4113/X sky130_fd_sc_hd__and2_1
XU$$4124 _555_/Q U$$4244/A2 U$$16/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4125/A sky130_fd_sc_hd__a22o_1
XFILLER_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4135 U$$4135/A U$$4197/B VGND VGND VPWR VPWR U$$4135/X sky130_fd_sc_hd__xor2_1
XU$$4146 _566_/Q U$$4244/A2 _567_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4147/A sky130_fd_sc_hd__a22o_1
XU$$3401 U$$3401/A U$$3403/B VGND VGND VPWR VPWR U$$3401/X sky130_fd_sc_hd__xor2_1
XU$$3412 U$$4508/A1 U$$3412/A2 _611_/Q U$$3412/B2 VGND VGND VPWR VPWR U$$3413/A sky130_fd_sc_hd__a22o_1
XFILLER_93_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4157 U$$4157/A U$$4197/B VGND VGND VPWR VPWR U$$4157/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_2 dadda_fa_4_113_2/A dadda_fa_4_113_2/B dadda_fa_4_113_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_114_0/CIN dadda_fa_5_113_1/CIN sky130_fd_sc_hd__fa_1
XU$$3423 U$$3423/A _665_/Q VGND VGND VPWR VPWR U$$3423/X sky130_fd_sc_hd__xor2_1
XU$$4168 _577_/Q U$$4198/A2 U$$4170/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4169/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4179 U$$4179/A U$$4197/B VGND VGND VPWR VPWR U$$4179/X sky130_fd_sc_hd__xor2_1
XU$$3434 U$$3434/A U$$3496/B VGND VGND VPWR VPWR U$$3434/X sky130_fd_sc_hd__xor2_1
XU$$2700 U$$2700/A _655_/Q VGND VGND VPWR VPWR U$$2700/X sky130_fd_sc_hd__xor2_1
XFILLER_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3445 U$$20/A1 U$$3429/X U$$979/B1 U$$3430/X VGND VGND VPWR VPWR U$$3446/A sky130_fd_sc_hd__a22o_1
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2711 U$$930/A1 U$$2607/X U$$932/A1 U$$2608/X VGND VGND VPWR VPWR U$$2712/A sky130_fd_sc_hd__a22o_1
XU$$3456 U$$3456/A U$$3496/B VGND VGND VPWR VPWR U$$3456/X sky130_fd_sc_hd__xor2_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_106_1 dadda_fa_4_106_1/A dadda_fa_4_106_1/B dadda_fa_4_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/B dadda_fa_5_106_1/B sky130_fd_sc_hd__fa_1
XU$$2722 U$$2722/A _655_/Q VGND VGND VPWR VPWR U$$2722/X sky130_fd_sc_hd__xor2_1
XU$$3467 U$$4289/A1 U$$3525/A2 U$$4289/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3468/A
+ sky130_fd_sc_hd__a22o_1
XU$$3478 U$$3478/A U$$3496/B VGND VGND VPWR VPWR U$$3478/X sky130_fd_sc_hd__xor2_1
XU$$2733 U$$4514/A1 U$$2607/X U$$4379/A1 U$$2608/X VGND VGND VPWR VPWR U$$2734/A sky130_fd_sc_hd__a22o_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2744 U$$2742/Y _656_/Q _655_/Q U$$2743/X U$$2740/Y VGND VGND VPWR VPWR U$$2744/X
+ sky130_fd_sc_hd__a32o_4
XU$$3489 U$$3900/A1 U$$3545/A2 U$$3489/B1 U$$3545/B2 VGND VGND VPWR VPWR U$$3490/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2755 U$$2755/A U$$2797/B VGND VGND VPWR VPWR U$$2755/X sky130_fd_sc_hd__xor2_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2766 U$$4273/A1 U$$2796/A2 U$$28/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2767/A sky130_fd_sc_hd__a22o_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2777 U$$2777/A U$$2797/B VGND VGND VPWR VPWR U$$2777/X sky130_fd_sc_hd__xor2_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2788 U$$4156/B1 U$$2868/A2 _573_/Q U$$2826/B2 VGND VGND VPWR VPWR U$$2789/A sky130_fd_sc_hd__a22o_1
XFILLER_18_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2799 U$$2799/A U$$2839/B VGND VGND VPWR VPWR U$$2799/X sky130_fd_sc_hd__xor2_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_127_0 dadda_fa_7_127_0/A dadda_fa_7_127_0/B dadda_fa_7_127_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_127_0/COUT _423_/D sky130_fd_sc_hd__fa_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_72_0 dadda_fa_2_72_0/A dadda_fa_2_72_0/B dadda_fa_2_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/B dadda_fa_3_72_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$706 final_adder.U$$706/A final_adder.U$$706/B VGND VGND VPWR VPWR
+ _252_/D sky130_fd_sc_hd__xor2_1
XFILLER_57_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$717 final_adder.U$$717/A final_adder.U$$717/B VGND VGND VPWR VPWR
+ _263_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$728 final_adder.U$$728/A final_adder.U$$728/B VGND VGND VPWR VPWR
+ _274_/D sky130_fd_sc_hd__xor2_1
XFILLER_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$739 final_adder.U$$739/A final_adder.U$$739/B VGND VGND VPWR VPWR
+ _285_/D sky130_fd_sc_hd__xor2_1
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3990 U$$3990/A U$$4044/B VGND VGND VPWR VPWR U$$3990/X sky130_fd_sc_hd__xor2_1
XFILLER_169_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR _560_/CLK sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_4_94_1 dadda_fa_4_94_1/A dadda_fa_4_94_1/B dadda_fa_4_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/B dadda_fa_5_94_1/B sky130_fd_sc_hd__fa_2
XFILLER_181_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_71_0 dadda_fa_7_71_0/A dadda_fa_7_71_0/B dadda_fa_7_71_0/CIN VGND VGND
+ VPWR VPWR _496_/D _367_/D sky130_fd_sc_hd__fa_2
XFILLER_118_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_87_0 dadda_fa_4_87_0/A dadda_fa_4_87_0/B dadda_fa_4_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/A dadda_fa_5_87_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_108_3 U$$4479/X input138/X dadda_fa_3_108_3/CIN VGND VGND VPWR VPWR dadda_fa_4_109_1/B
+ dadda_fa_4_108_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_133_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput270 _279_/Q VGND VGND VPWR VPWR o[111] sky130_fd_sc_hd__buf_2
Xoutput281 _289_/Q VGND VGND VPWR VPWR o[121] sky130_fd_sc_hd__buf_2
XFILLER_58_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput292 _184_/Q VGND VGND VPWR VPWR o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2007 U$$2007/A U$$2055/A VGND VGND VPWR VPWR U$$2007/X sky130_fd_sc_hd__xor2_1
XFILLER_28_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2018 U$$785/A1 U$$2048/A2 U$$924/A1 U$$2048/B2 VGND VGND VPWR VPWR U$$2019/A sky130_fd_sc_hd__a22o_1
XU$$2029 U$$2029/A U$$2055/A VGND VGND VPWR VPWR U$$2029/X sky130_fd_sc_hd__xor2_1
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1306 U$$1306/A U$$1369/A VGND VGND VPWR VPWR U$$1306/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1317 U$$84/A1 U$$1367/A2 U$$908/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1318/A sky130_fd_sc_hd__a22o_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1328 U$$1328/A U$$1342/B VGND VGND VPWR VPWR U$$1328/X sky130_fd_sc_hd__xor2_1
XU$$1339 U$$928/A1 U$$1367/A2 _602_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1340/A sky130_fd_sc_hd__a22o_1
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_205_ _448_/CLK _205_/D VGND VGND VPWR VPWR _205_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_51_5 dadda_fa_2_51_5/A dadda_fa_2_51_5/B dadda_fa_2_51_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_2/A dadda_fa_4_51_0/A sky130_fd_sc_hd__fa_2
X_762__814 VGND VGND VPWR VPWR _762__814/HI U$$4116/A1 sky130_fd_sc_hd__conb_1
XFILLER_94_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_44_4 dadda_fa_2_44_4/A dadda_fa_2_44_4/B dadda_fa_2_44_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/CIN dadda_fa_3_44_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3220 U$$3220/A U$$3244/B VGND VGND VPWR VPWR U$$3220/X sky130_fd_sc_hd__xor2_1
XFILLER_19_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3231 _588_/Q U$$3155/X _589_/Q U$$3156/X VGND VGND VPWR VPWR U$$3232/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_6_3_0 U$$13/X U$$146/X VGND VGND VPWR VPWR dadda_fa_7_4_0/B dadda_ha_6_3_0/SUM
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$13 _437_/Q _309_/Q VGND VGND VPWR VPWR final_adder.U$$141/B1 final_adder.U$$635/A
+ sky130_fd_sc_hd__ha_1
XFILLER_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3242 U$$3242/A _663_/Q VGND VGND VPWR VPWR U$$3242/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$24 _448_/Q _320_/Q VGND VGND VPWR VPWR final_adder.U$$519/B1 final_adder.U$$646/A
+ sky130_fd_sc_hd__ha_1
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3253 U$$4486/A1 U$$3155/X U$$787/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3254/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$35 _459_/Q _331_/Q VGND VGND VPWR VPWR final_adder.U$$163/B1 final_adder.U$$657/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_37_3 U$$1943/X U$$2076/X U$$2209/X VGND VGND VPWR VPWR dadda_fa_3_38_1/B
+ dadda_fa_3_37_3/B sky130_fd_sc_hd__fa_1
XU$$3264 U$$3264/A U$$3270/B VGND VGND VPWR VPWR U$$3264/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$46 _470_/Q _342_/Q VGND VGND VPWR VPWR final_adder.U$$541/B1 final_adder.U$$668/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$57 _481_/Q _353_/Q VGND VGND VPWR VPWR final_adder.U$$185/B1 final_adder.U$$679/A
+ sky130_fd_sc_hd__ha_1
XU$$3275 U$$4508/A1 U$$3155/X _611_/Q U$$3156/X VGND VGND VPWR VPWR U$$3276/A sky130_fd_sc_hd__a22o_1
XU$$2530 U$$64/A1 U$$2574/A2 U$$66/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2531/A sky130_fd_sc_hd__a22o_1
XU$$2541 U$$2541/A U$$2585/B VGND VGND VPWR VPWR U$$2541/X sky130_fd_sc_hd__xor2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_803__855 VGND VGND VPWR VPWR _803__855/HI U$$4451/B sky130_fd_sc_hd__conb_1
XU$$3286 U$$3286/A _663_/Q VGND VGND VPWR VPWR U$$3286/X sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$68 _492_/Q _364_/Q VGND VGND VPWR VPWR final_adder.U$$563/B1 final_adder.U$$690/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3297 U$$3297/A U$$3413/B VGND VGND VPWR VPWR U$$3297/X sky130_fd_sc_hd__xor2_1
XU$$2552 U$$86/A1 U$$2584/A2 U$$88/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2553/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$79 _503_/Q _375_/Q VGND VGND VPWR VPWR final_adder.U$$207/B1 final_adder.U$$701/A
+ sky130_fd_sc_hd__ha_1
XU$$2563 U$$2563/A U$$2585/B VGND VGND VPWR VPWR U$$2563/X sky130_fd_sc_hd__xor2_1
XU$$2574 U$$930/A1 U$$2574/A2 U$$932/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2575/A sky130_fd_sc_hd__a22o_1
XU$$1840 U$$1840/A U$$1856/B VGND VGND VPWR VPWR U$$1840/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2585 U$$2585/A U$$2585/B VGND VGND VPWR VPWR U$$2585/X sky130_fd_sc_hd__xor2_1
XU$$1851 U$$892/A1 U$$1903/A2 U$$892/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1852/A sky130_fd_sc_hd__a22o_1
XU$$2596 U$$4514/A1 U$$2470/X U$$4379/A1 U$$2471/X VGND VGND VPWR VPWR U$$2597/A sky130_fd_sc_hd__a22o_1
XU$$1862 U$$1862/A U$$1918/A VGND VGND VPWR VPWR U$$1862/X sky130_fd_sc_hd__xor2_1
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1873 U$$4476/A1 U$$1785/X U$$94/A1 U$$1786/X VGND VGND VPWR VPWR U$$1874/A sky130_fd_sc_hd__a22o_1
XU$$1884 U$$1884/A U$$1904/B VGND VGND VPWR VPWR U$$1884/X sky130_fd_sc_hd__xor2_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1895 U$$936/A1 U$$1785/X _606_/Q U$$1786/X VGND VGND VPWR VPWR U$$1896/A sky130_fd_sc_hd__a22o_1
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$503 final_adder.U$$8/SUM final_adder.U$$630/B final_adder.U$$8/COUT
+ VGND VGND VPWR VPWR final_adder.U$$631/B sky130_fd_sc_hd__a21o_1
XFILLER_57_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$525 final_adder.U$$652/A final_adder.U$$652/B final_adder.U$$525/B1
+ VGND VGND VPWR VPWR final_adder.U$$653/B sky130_fd_sc_hd__a21o_1
XFILLER_57_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater740 _561_/Q VGND VGND VPWR VPWR U$$4273/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$547 final_adder.U$$674/A final_adder.U$$674/B final_adder.U$$547/B1
+ VGND VGND VPWR VPWR final_adder.U$$675/B sky130_fd_sc_hd__a21o_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater751 _556_/Q VGND VGND VPWR VPWR U$$14/B1 sky130_fd_sc_hd__buf_12
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$569 final_adder.U$$696/A final_adder.U$$696/B final_adder.U$$569/B1
+ VGND VGND VPWR VPWR final_adder.U$$697/B sky130_fd_sc_hd__a21o_1
XU$$408 U$$819/A1 U$$278/X U$$408/B1 U$$279/X VGND VGND VPWR VPWR U$$409/A sky130_fd_sc_hd__a22o_1
XU$$419 _552_/Q U$$491/A2 U$$969/A1 U$$416/X VGND VGND VPWR VPWR U$$420/A sky130_fd_sc_hd__a22o_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_113_1 U$$3824/X U$$3957/X U$$4090/X VGND VGND VPWR VPWR dadda_fa_4_114_2/A
+ dadda_fa_4_113_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_0 U$$3544/X U$$3677/X U$$3810/X VGND VGND VPWR VPWR dadda_fa_4_107_0/B
+ dadda_fa_4_106_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_54_3 dadda_fa_3_54_3/A dadda_fa_3_54_3/B dadda_fa_3_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/B dadda_fa_4_54_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_134_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_47_2 dadda_fa_3_47_2/A dadda_fa_3_47_2/B dadda_fa_3_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/A dadda_fa_4_47_2/B sky130_fd_sc_hd__fa_1
XFILLER_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$920 U$$98/A1 U$$826/X U$$98/B1 U$$827/X VGND VGND VPWR VPWR U$$921/A sky130_fd_sc_hd__a22o_1
XU$$931 U$$931/A U$$943/B VGND VGND VPWR VPWR U$$931/X sky130_fd_sc_hd__xor2_1
XU$$942 U$$942/A1 U$$826/X U$$944/A1 U$$827/X VGND VGND VPWR VPWR U$$943/A sky130_fd_sc_hd__a22o_1
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_17_0 dadda_fa_6_17_0/A dadda_fa_6_17_0/B dadda_fa_6_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_18_0/B dadda_fa_7_17_0/CIN sky130_fd_sc_hd__fa_1
XU$$953 U$$953/A _629_/Q VGND VGND VPWR VPWR U$$953/X sky130_fd_sc_hd__xor2_1
XFILLER_91_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1103 U$$1103/A U$$1189/B VGND VGND VPWR VPWR U$$1103/X sky130_fd_sc_hd__xor2_1
XU$$964 U$$962/B U$$959/A _630_/Q U$$959/Y VGND VGND VPWR VPWR U$$964/X sky130_fd_sc_hd__a22o_4
XFILLER_44_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1114 U$$18/A1 U$$1200/A2 U$$20/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1115/A sky130_fd_sc_hd__a22o_1
XU$$975 U$$16/A1 U$$999/A2 U$$975/B1 U$$999/B2 VGND VGND VPWR VPWR U$$976/A sky130_fd_sc_hd__a22o_1
XU$$1125 U$$1125/A U$$1189/B VGND VGND VPWR VPWR U$$1125/X sky130_fd_sc_hd__xor2_1
XU$$986 U$$986/A U$$992/B VGND VGND VPWR VPWR U$$986/X sky130_fd_sc_hd__xor2_1
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$997 U$$38/A1 U$$963/X U$$40/A1 U$$999/B2 VGND VGND VPWR VPWR U$$998/A sky130_fd_sc_hd__a22o_1
XU$$1136 U$$3191/A1 U$$1200/A2 U$$3876/B1 U$$1200/B2 VGND VGND VPWR VPWR U$$1137/A
+ sky130_fd_sc_hd__a22o_1
XU$$1147 U$$1147/A U$$1167/B VGND VGND VPWR VPWR U$$1147/X sky130_fd_sc_hd__xor2_1
XU$$1158 U$$3624/A1 U$$1218/A2 U$$3900/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1159/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1169 U$$1169/A U$$1232/A VGND VGND VPWR VPWR U$$1169/X sky130_fd_sc_hd__xor2_1
XFILLER_129_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_42_1 U$$2352/X U$$2485/X U$$2618/X VGND VGND VPWR VPWR dadda_fa_3_43_0/CIN
+ dadda_fa_3_42_2/CIN sky130_fd_sc_hd__fa_1
XU$$3050 U$$4283/A1 U$$3090/A2 U$$4285/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3051/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3061 U$$3061/A U$$3129/B VGND VGND VPWR VPWR U$$3061/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_0 U$$343/X U$$476/X U$$609/X VGND VGND VPWR VPWR dadda_fa_3_36_0/B
+ dadda_fa_3_35_2/B sky130_fd_sc_hd__fa_2
XU$$3072 U$$4442/A1 U$$3090/A2 U$$4170/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3073/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3083 U$$3083/A U$$3109/B VGND VGND VPWR VPWR U$$3083/X sky130_fd_sc_hd__xor2_1
XU$$3094 U$$902/A1 U$$3146/A2 U$$902/B1 U$$3146/B2 VGND VGND VPWR VPWR U$$3095/A sky130_fd_sc_hd__a22o_1
XU$$2360 U$$2360/A U$$2432/B VGND VGND VPWR VPWR U$$2360/X sky130_fd_sc_hd__xor2_1
XU$$2371 U$$4289/A1 U$$2421/A2 U$$4289/B1 U$$2421/B2 VGND VGND VPWR VPWR U$$2372/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2382 U$$2382/A U$$2436/B VGND VGND VPWR VPWR U$$2382/X sky130_fd_sc_hd__xor2_1
XFILLER_22_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2393 U$$3900/A1 U$$2421/A2 U$$3489/B1 U$$2421/B2 VGND VGND VPWR VPWR U$$2394/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1670 U$$4273/A1 U$$1726/A2 U$$987/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1671/A
+ sky130_fd_sc_hd__a22o_1
XU$$1681 U$$1681/A U$$1727/B VGND VGND VPWR VPWR U$$1681/X sky130_fd_sc_hd__xor2_1
XFILLER_10_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1692 U$$48/A1 U$$1726/A2 U$$50/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1693/A sky130_fd_sc_hd__a22o_1
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_87_3 U$$2841/X U$$2974/X U$$3107/X VGND VGND VPWR VPWR dadda_fa_2_88_4/A
+ dadda_fa_2_87_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_64_2 dadda_fa_4_64_2/A dadda_fa_4_64_2/B dadda_fa_4_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/CIN dadda_fa_5_64_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_57_1 dadda_fa_4_57_1/A dadda_fa_4_57_1/B dadda_fa_4_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/B dadda_fa_5_57_1/B sky130_fd_sc_hd__fa_1
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$300 final_adder.U$$300/A final_adder.U$$300/B VGND VGND VPWR VPWR
+ final_adder.U$$342/B sky130_fd_sc_hd__and2_1
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$311 final_adder.U$$310/A final_adder.U$$237/X final_adder.U$$239/X
+ VGND VGND VPWR VPWR final_adder.U$$311/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_34_0 dadda_fa_7_34_0/A dadda_fa_7_34_0/B dadda_fa_7_34_0/CIN VGND VGND
+ VPWR VPWR _459_/D _330_/D sky130_fd_sc_hd__fa_2
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$322 final_adder.U$$322/A final_adder.U$$322/B VGND VGND VPWR VPWR
+ final_adder.U$$322/X sky130_fd_sc_hd__and2_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$333 final_adder.U$$332/A final_adder.U$$281/X final_adder.U$$283/X
+ VGND VGND VPWR VPWR final_adder.U$$333/X sky130_fd_sc_hd__a21o_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$344 final_adder.U$$344/A final_adder.U$$344/B VGND VGND VPWR VPWR
+ final_adder.U$$364/B sky130_fd_sc_hd__and2_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$355 final_adder.U$$354/A final_adder.U$$325/X final_adder.U$$327/X
+ VGND VGND VPWR VPWR final_adder.U$$355/X sky130_fd_sc_hd__a21o_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater570 _645_/Q VGND VGND VPWR VPWR U$$2055/A sky130_fd_sc_hd__buf_12
XU$$205 U$$68/A1 U$$141/X U$$68/B1 U$$142/X VGND VGND VPWR VPWR U$$206/A sky130_fd_sc_hd__a22o_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$377 final_adder.U$$370/X final_adder.U$$654/B final_adder.U$$371/X
+ VGND VGND VPWR VPWR final_adder.U$$686/B sky130_fd_sc_hd__a21o_4
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$216 U$$216/A U$$274/A VGND VGND VPWR VPWR U$$216/X sky130_fd_sc_hd__xor2_1
Xrepeater581 U$$1479/B VGND VGND VPWR VPWR U$$1461/B sky130_fd_sc_hd__buf_12
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$227 U$$90/A1 U$$141/X U$$92/A1 U$$142/X VGND VGND VPWR VPWR U$$228/A sky130_fd_sc_hd__a22o_1
Xrepeater592 _631_/Q VGND VGND VPWR VPWR U$$998/B sky130_fd_sc_hd__buf_12
XFILLER_45_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$399 final_adder.U$$362/B final_adder.U$$702/B final_adder.U$$341/X
+ VGND VGND VPWR VPWR final_adder.U$$710/B sky130_fd_sc_hd__a21o_1
XU$$238 U$$238/A U$$274/A VGND VGND VPWR VPWR U$$238/X sky130_fd_sc_hd__xor2_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$249 U$$934/A1 U$$141/X U$$799/A1 U$$142/X VGND VGND VPWR VPWR U$$250/A sky130_fd_sc_hd__a22o_1
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_470_ _471_/CLK _470_/D VGND VGND VPWR VPWR _470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_75_1 U$$1221/X U$$1354/X U$$1487/X VGND VGND VPWR VPWR dadda_fa_1_76_8/B
+ dadda_fa_2_75_0/A sky130_fd_sc_hd__fa_2
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_52_0 dadda_fa_3_52_0/A dadda_fa_3_52_0/B dadda_fa_3_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/B dadda_fa_4_52_1/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_0_68_0 _680__900/HI U$$409/X U$$542/X VGND VGND VPWR VPWR dadda_fa_1_69_5/CIN
+ dadda_fa_1_68_7/B sky130_fd_sc_hd__fa_2
XFILLER_64_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$750 U$$750/A U$$778/B VGND VGND VPWR VPWR U$$750/X sky130_fd_sc_hd__xor2_1
X_668_ _679_/CLK _668_/D VGND VGND VPWR VPWR _668_/Q sky130_fd_sc_hd__dfxtp_1
XU$$761 U$$76/A1 U$$785/A2 U$$76/B1 U$$785/B2 VGND VGND VPWR VPWR U$$762/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$772 U$$772/A U$$822/A VGND VGND VPWR VPWR U$$772/X sky130_fd_sc_hd__xor2_1
XU$$783 U$$98/A1 U$$817/A2 U$$98/B1 U$$817/B2 VGND VGND VPWR VPWR U$$784/A sky130_fd_sc_hd__a22o_1
XFILLER_56_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$794 U$$794/A _627_/Q VGND VGND VPWR VPWR U$$794/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_599_ _601_/CLK _599_/D VGND VGND VPWR VPWR _599_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_clk _560_/CLK VGND VGND VPWR VPWR _679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_176_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_97_2 U$$3127/X U$$3260/X U$$3393/X VGND VGND VPWR VPWR dadda_fa_3_98_1/A
+ dadda_fa_3_97_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_74_1 dadda_fa_5_74_1/A dadda_fa_5_74_1/B dadda_fa_5_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/B dadda_fa_7_74_0/A sky130_fd_sc_hd__fa_1
XFILLER_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_67_0 dadda_fa_5_67_0/A dadda_fa_5_67_0/B dadda_fa_5_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/A dadda_fa_6_67_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_768__820 VGND VGND VPWR VPWR _768__820/HI U$$4386/A sky130_fd_sc_hd__conb_1
XFILLER_101_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_66_8 dadda_fa_1_66_8/A dadda_fa_1_66_8/B dadda_fa_1_66_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_3/A dadda_fa_3_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_6_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_809__861 VGND VGND VPWR VPWR _809__861/HI U$$4463/B sky130_fd_sc_hd__conb_1
XFILLER_6_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_59_7 dadda_fa_1_59_7/A dadda_fa_1_59_7/B dadda_fa_1_59_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_2/CIN dadda_fa_2_59_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_6_0 input223/X dadda_fa_6_6_0/B dadda_fa_6_6_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_7_7_0/B dadda_fa_7_6_0/CIN sky130_fd_sc_hd__fa_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2190 U$$2190/A U$$2192/A VGND VGND VPWR VPWR U$$2190/X sky130_fd_sc_hd__xor2_1
XFILLER_148_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_92_1 U$$2319/X U$$2452/X U$$2585/X VGND VGND VPWR VPWR dadda_fa_2_93_5/A
+ dadda_fa_2_92_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_85_0 U$$1506/Y U$$1640/X U$$1773/X VGND VGND VPWR VPWR dadda_fa_2_86_2/B
+ dadda_fa_2_85_4/B sky130_fd_sc_hd__fa_1
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4509 U$$4509/A U$$4509/B VGND VGND VPWR VPWR U$$4509/X sky130_fd_sc_hd__xor2_2
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$130 final_adder.U$$625/A final_adder.U$$624/A VGND VGND VPWR VPWR
+ final_adder.U$$130/X sky130_fd_sc_hd__and2_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3808 U$$3808/A U$$3835/A VGND VGND VPWR VPWR U$$3808/X sky130_fd_sc_hd__xor2_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$141 final_adder.U$$635/A final_adder.U$$507/B1 final_adder.U$$141/B1
+ VGND VGND VPWR VPWR final_adder.U$$141/X sky130_fd_sc_hd__a21o_1
XFILLER_18_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3819 U$$4504/A1 U$$3703/X U$$4506/A1 U$$3704/X VGND VGND VPWR VPWR U$$3820/A sky130_fd_sc_hd__a22o_1
XFILLER_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$152 final_adder.U$$647/A final_adder.U$$646/A VGND VGND VPWR VPWR
+ final_adder.U$$268/B sky130_fd_sc_hd__and2_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$163 final_adder.U$$657/A final_adder.U$$529/B1 final_adder.U$$163/B1
+ VGND VGND VPWR VPWR final_adder.U$$163/X sky130_fd_sc_hd__a21o_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$174 final_adder.U$$669/A final_adder.U$$668/A VGND VGND VPWR VPWR
+ final_adder.U$$278/A sky130_fd_sc_hd__and2_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$185 final_adder.U$$679/A final_adder.U$$551/B1 final_adder.U$$185/B1
+ VGND VGND VPWR VPWR final_adder.U$$185/X sky130_fd_sc_hd__a21o_1
XFILLER_166_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$196 final_adder.U$$691/A final_adder.U$$690/A VGND VGND VPWR VPWR
+ final_adder.U$$290/B sky130_fd_sc_hd__and2_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_522_ _537_/CLK _522_/D VGND VGND VPWR VPWR _522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_126_0 _709__929/HI U$$4382/X VGND VGND VPWR VPWR dadda_fa_7_127_0/A dadda_fa_7_126_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ _462_/CLK _453_/D VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _535_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_384_ _387_/CLK _384_/D VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_84_0 dadda_fa_6_84_0/A dadda_fa_6_84_0/B dadda_fa_6_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_85_0/B dadda_fa_7_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_182_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput170 c[21] VGND VGND VPWR VPWR input170/X sky130_fd_sc_hd__buf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput181 c[31] VGND VGND VPWR VPWR input181/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput192 c[41] VGND VGND VPWR VPWR input192/X sky130_fd_sc_hd__buf_2
XFILLER_37_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$580 U$$32/A1 U$$682/A2 U$$34/A1 U$$553/X VGND VGND VPWR VPWR U$$581/A sky130_fd_sc_hd__a22o_1
XU$$591 U$$591/A U$$623/B VGND VGND VPWR VPWR U$$591/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_43_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _527_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_71_6 input225/X dadda_fa_1_71_6/B dadda_fa_1_71_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_72_2/B dadda_fa_2_71_5/B sky130_fd_sc_hd__fa_1
XFILLER_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_64_5 input217/X dadda_fa_1_64_5/B dadda_fa_1_64_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_65_2/A dadda_fa_2_64_5/A sky130_fd_sc_hd__fa_2
XFILLER_74_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_4 U$$2781/X U$$2914/X U$$3047/X VGND VGND VPWR VPWR dadda_fa_2_58_1/CIN
+ dadda_fa_2_57_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_27_2 dadda_fa_4_27_2/A dadda_fa_4_27_2/B dadda_fa_4_27_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/CIN dadda_fa_5_27_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _509_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4306 U$$4306/A U$$4384/A VGND VGND VPWR VPWR U$$4306/X sky130_fd_sc_hd__xor2_1
XU$$4317 U$$70/A1 U$$4377/A2 U$$70/B1 U$$4377/B2 VGND VGND VPWR VPWR U$$4318/A sky130_fd_sc_hd__a22o_1
XFILLER_120_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4328 U$$4328/A U$$4332/B VGND VGND VPWR VPWR U$$4328/X sky130_fd_sc_hd__xor2_1
XU$$4339 U$$4476/A1 U$$4381/A2 U$$94/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4340/A sky130_fd_sc_hd__a22o_1
XFILLER_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3605 U$$3605/A U$$3625/B VGND VGND VPWR VPWR U$$3605/X sky130_fd_sc_hd__xor2_1
XU$$3616 U$$4438/A1 U$$3678/A2 _576_/Q U$$3678/B2 VGND VGND VPWR VPWR U$$3617/A sky130_fd_sc_hd__a22o_1
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3627 U$$3627/A _669_/Q VGND VGND VPWR VPWR U$$3627/X sky130_fd_sc_hd__xor2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3638 U$$76/A1 U$$3668/A2 _587_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3639/A sky130_fd_sc_hd__a22o_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2904 U$$2904/A U$$2960/B VGND VGND VPWR VPWR U$$2904/X sky130_fd_sc_hd__xor2_1
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3649 U$$3649/A U$$3699/A VGND VGND VPWR VPWR U$$3649/X sky130_fd_sc_hd__xor2_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2915 U$$4285/A1 U$$2975/A2 U$$4424/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2916/A
+ sky130_fd_sc_hd__a22o_1
XU$$2926 U$$2926/A U$$2996/B VGND VGND VPWR VPWR U$$2926/X sky130_fd_sc_hd__xor2_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2937 _578_/Q U$$2975/A2 U$$3624/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2938/A sky130_fd_sc_hd__a22o_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2948 U$$2948/A U$$3004/B VGND VGND VPWR VPWR U$$2948/X sky130_fd_sc_hd__xor2_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ _509_/CLK _505_/D VGND VGND VPWR VPWR _505_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_3_22_1 U$$716/X U$$849/X U$$982/X VGND VGND VPWR VPWR dadda_fa_4_23_0/CIN
+ dadda_fa_4_22_2/A sky130_fd_sc_hd__fa_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2959 U$$902/B1 U$$2975/A2 U$$84/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2960/A sky130_fd_sc_hd__a22o_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk _369_/CLK VGND VGND VPWR VPWR _480_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_436_ _455_/CLK _436_/D VGND VGND VPWR VPWR _436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_367_ _367_/CLK _367_/D VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_298_ _429_/CLK _298_/D VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_81_5 dadda_fa_2_81_5/A dadda_fa_2_81_5/B dadda_fa_2_81_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_2/A dadda_fa_4_81_0/A sky130_fd_sc_hd__fa_1
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_4 dadda_fa_2_74_4/A dadda_fa_2_74_4/B dadda_fa_2_74_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/CIN dadda_fa_3_74_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_730__782 VGND VGND VPWR VPWR _730__782/HI U$$2198/A1 sky130_fd_sc_hd__conb_1
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_67_3 dadda_fa_2_67_3/A dadda_fa_2_67_3/B dadda_fa_2_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/B dadda_fa_3_67_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_37_1 dadda_fa_5_37_1/A dadda_fa_5_37_1/B dadda_fa_5_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/B dadda_fa_7_37_0/A sky130_fd_sc_hd__fa_2
XFILLER_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_16_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _458_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_111_1 dadda_fa_5_111_1/A dadda_fa_5_111_1/B dadda_fa_5_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/B dadda_fa_7_111_0/A sky130_fd_sc_hd__fa_2
XFILLER_34_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_104_0 dadda_fa_5_104_0/A dadda_fa_5_104_0/B dadda_fa_5_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/A dadda_fa_6_104_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_2 U$$3190/X U$$3323/X U$$3456/X VGND VGND VPWR VPWR dadda_fa_2_63_1/A
+ dadda_fa_2_62_4/A sky130_fd_sc_hd__fa_2
XFILLER_102_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_55_1 U$$1181/X U$$1314/X U$$1447/X VGND VGND VPWR VPWR dadda_fa_2_56_0/CIN
+ dadda_fa_2_55_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_32_0 dadda_fa_4_32_0/A dadda_fa_4_32_0/B dadda_fa_4_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/A dadda_fa_5_32_1/A sky130_fd_sc_hd__fa_1
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_48_0 U$$103/X U$$236/X U$$369/X VGND VGND VPWR VPWR dadda_fa_2_49_1/A
+ dadda_fa_2_48_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_103_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_221_ _474_/CLK _221_/D VGND VGND VPWR VPWR _221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_84_3 dadda_fa_3_84_3/A dadda_fa_3_84_3/B dadda_fa_3_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/B dadda_fa_4_84_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_714__766 VGND VGND VPWR VPWR _714__766/HI U$$1239/A1 sky130_fd_sc_hd__conb_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_77_2 dadda_fa_3_77_2/A dadda_fa_3_77_2/B dadda_fa_3_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/A dadda_fa_4_77_2/B sky130_fd_sc_hd__fa_2
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_47_0 dadda_fa_6_47_0/A dadda_fa_6_47_0/B dadda_fa_6_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_48_0/B dadda_fa_7_47_0/CIN sky130_fd_sc_hd__fa_1
XU$$4103 _613_/Q U$$4107/A2 U$$4379/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4104/A sky130_fd_sc_hd__a22o_1
XU$$4114 U$$4112/Y _676_/Q _675_/Q U$$4113/X U$$4110/Y VGND VGND VPWR VPWR U$$4114/X
+ sky130_fd_sc_hd__a32o_4
XU$$4125 U$$4125/A _677_/Q VGND VGND VPWR VPWR U$$4125/X sky130_fd_sc_hd__xor2_1
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4136 U$$4273/A1 U$$4114/X _562_/Q U$$4198/B2 VGND VGND VPWR VPWR U$$4137/A sky130_fd_sc_hd__a22o_1
XU$$4147 U$$4147/A U$$4246/A VGND VGND VPWR VPWR U$$4147/X sky130_fd_sc_hd__xor2_1
XFILLER_59_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3402 _605_/Q U$$3292/X U$$4500/A1 U$$3293/X VGND VGND VPWR VPWR U$$3403/A sky130_fd_sc_hd__a22o_1
XU$$3413 U$$3413/A U$$3413/B VGND VGND VPWR VPWR U$$3413/X sky130_fd_sc_hd__xor2_1
XU$$4158 _572_/Q U$$4198/A2 U$$735/A1 U$$4198/B2 VGND VGND VPWR VPWR U$$4159/A sky130_fd_sc_hd__a22o_1
XU$$3424 _665_/Q VGND VGND VPWR VPWR U$$3424/Y sky130_fd_sc_hd__inv_1
XFILLER_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4169 U$$4169/A U$$4247/A VGND VGND VPWR VPWR U$$4169/X sky130_fd_sc_hd__xor2_1
XU$$3435 _553_/Q U$$3525/A2 U$$4122/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3436/A sky130_fd_sc_hd__a22o_1
XU$$2701 _597_/Q U$$2607/X _598_/Q U$$2608/X VGND VGND VPWR VPWR U$$2702/A sky130_fd_sc_hd__a22o_1
XU$$3446 U$$3446/A U$$3561/A VGND VGND VPWR VPWR U$$3446/X sky130_fd_sc_hd__xor2_1
XFILLER_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2712 U$$2712/A _655_/Q VGND VGND VPWR VPWR U$$2712/X sky130_fd_sc_hd__xor2_1
XU$$3457 U$$30/B1 U$$3525/A2 U$$3457/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3458/A sky130_fd_sc_hd__a22o_1
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2723 _608_/Q U$$2607/X _609_/Q U$$2608/X VGND VGND VPWR VPWR U$$2724/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_2 dadda_fa_4_106_2/A dadda_fa_4_106_2/B dadda_fa_4_106_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/CIN dadda_fa_5_106_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3468 U$$3468/A U$$3496/B VGND VGND VPWR VPWR U$$3468/X sky130_fd_sc_hd__xor2_1
XU$$3479 _575_/Q U$$3545/A2 U$$4303/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3480/A sky130_fd_sc_hd__a22o_1
XU$$2734 U$$2734/A _655_/Q VGND VGND VPWR VPWR U$$2734/X sky130_fd_sc_hd__xor2_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2745 U$$2743/B _655_/Q _656_/Q U$$2740/Y VGND VGND VPWR VPWR U$$2745/X sky130_fd_sc_hd__a22o_4
XU$$2756 _556_/Q U$$2796/A2 U$$4265/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2757/A sky130_fd_sc_hd__a22o_1
XFILLER_34_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2767 U$$2767/A U$$2797/B VGND VGND VPWR VPWR U$$2767/X sky130_fd_sc_hd__xor2_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2778 U$$4285/A1 U$$2796/A2 U$$3191/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2779/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2789 U$$2789/A U$$2839/B VGND VGND VPWR VPWR U$$2789/X sky130_fd_sc_hd__xor2_1
XFILLER_18_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_419_ _615_/CLK _419_/D VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_5_clk _369_/CLK VGND VGND VPWR VPWR _469_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_72_1 dadda_fa_2_72_1/A dadda_fa_2_72_1/B dadda_fa_2_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/CIN dadda_fa_3_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_25_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_65_0 dadda_fa_2_65_0/A dadda_fa_2_65_0/B dadda_fa_2_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/B dadda_fa_3_65_2/B sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$707 final_adder.U$$707/A final_adder.U$$707/B VGND VGND VPWR VPWR
+ _253_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$718 final_adder.U$$718/A final_adder.U$$718/B VGND VGND VPWR VPWR
+ _264_/D sky130_fd_sc_hd__xor2_1
XFILLER_57_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$729 final_adder.U$$729/A final_adder.U$$729/B VGND VGND VPWR VPWR
+ _275_/D sky130_fd_sc_hd__xor2_1
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_704__924 VGND VGND VPWR VPWR _704__924/HI _704__924/LO sky130_fd_sc_hd__conb_1
XFILLER_80_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3980 U$$3980/A U$$4044/B VGND VGND VPWR VPWR U$$3980/X sky130_fd_sc_hd__xor2_1
XU$$3991 _557_/Q U$$4045/A2 U$$842/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$3992/A sky130_fd_sc_hd__a22o_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_94_2 dadda_fa_4_94_2/A dadda_fa_4_94_2/B dadda_fa_4_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/CIN dadda_fa_5_94_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_192_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_87_1 dadda_fa_4_87_1/A dadda_fa_4_87_1/B dadda_fa_4_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/B dadda_fa_5_87_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_64_0 dadda_fa_7_64_0/A dadda_fa_7_64_0/B dadda_fa_7_64_0/CIN VGND VGND
+ VPWR VPWR _489_/D _360_/D sky130_fd_sc_hd__fa_2
XFILLER_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput260 _270_/Q VGND VGND VPWR VPWR o[102] sky130_fd_sc_hd__buf_2
XFILLER_161_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput271 _280_/Q VGND VGND VPWR VPWR o[112] sky130_fd_sc_hd__buf_2
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput282 _290_/Q VGND VGND VPWR VPWR o[122] sky130_fd_sc_hd__buf_2
Xoutput293 _185_/Q VGND VGND VPWR VPWR o[17] sky130_fd_sc_hd__buf_2
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2008 U$$912/A1 U$$2036/A2 U$$914/A1 U$$2036/B2 VGND VGND VPWR VPWR U$$2009/A sky130_fd_sc_hd__a22o_1
XU$$2019 U$$2019/A U$$2055/A VGND VGND VPWR VPWR U$$2019/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1307 U$$74/A1 U$$1341/A2 U$$2953/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1308/A sky130_fd_sc_hd__a22o_1
XU$$1318 U$$1318/A U$$1369/A VGND VGND VPWR VPWR U$$1318/X sky130_fd_sc_hd__xor2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1329 U$$94/B1 U$$1341/A2 U$$98/A1 U$$1341/B2 VGND VGND VPWR VPWR U$$1330/A sky130_fd_sc_hd__a22o_1
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_204_ _448_/CLK _204_/D VGND VGND VPWR VPWR _204_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_82_0 dadda_fa_3_82_0/A dadda_fa_3_82_0/B dadda_fa_3_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/B dadda_fa_4_82_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_174_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3210 U$$3210/A U$$3244/B VGND VGND VPWR VPWR U$$3210/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3221 _583_/Q U$$3243/A2 _584_/Q U$$3243/B2 VGND VGND VPWR VPWR U$$3222/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_111_0 U$$4485/X input142/X dadda_fa_4_111_0/CIN VGND VGND VPWR VPWR dadda_fa_5_112_0/A
+ dadda_fa_5_111_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_44_5 dadda_fa_2_44_5/A dadda_fa_2_44_5/B dadda_fa_2_44_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_2/A dadda_fa_4_44_0/A sky130_fd_sc_hd__fa_2
XU$$3232 U$$3232/A U$$3270/B VGND VGND VPWR VPWR U$$3232/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$14 _438_/Q _310_/Q VGND VGND VPWR VPWR final_adder.U$$509/B1 final_adder.U$$636/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$25 _449_/Q _321_/Q VGND VGND VPWR VPWR final_adder.U$$153/B1 final_adder.U$$647/A
+ sky130_fd_sc_hd__ha_1
XFILLER_47_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3243 U$$4476/A1 U$$3243/A2 _595_/Q U$$3243/B2 VGND VGND VPWR VPWR U$$3244/A sky130_fd_sc_hd__a22o_1
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3254 U$$3254/A _663_/Q VGND VGND VPWR VPWR U$$3254/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$36 _460_/Q _332_/Q VGND VGND VPWR VPWR final_adder.U$$531/B1 final_adder.U$$658/A
+ sky130_fd_sc_hd__ha_1
XFILLER_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_37_4 U$$2342/X U$$2475/X input187/X VGND VGND VPWR VPWR dadda_fa_3_38_1/CIN
+ dadda_fa_3_37_3/CIN sky130_fd_sc_hd__fa_1
XU$$3265 _605_/Q U$$3155/X U$$4500/A1 U$$3156/X VGND VGND VPWR VPWR U$$3266/A sky130_fd_sc_hd__a22o_1
XFILLER_111_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2520 U$$876/A1 U$$2534/A2 U$$878/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2521/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$47 _471_/Q _343_/Q VGND VGND VPWR VPWR final_adder.U$$175/B1 final_adder.U$$669/A
+ sky130_fd_sc_hd__ha_1
X_842__894 VGND VGND VPWR VPWR _842__894/HI U$$691/A1 sky130_fd_sc_hd__conb_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3276 U$$3276/A _663_/Q VGND VGND VPWR VPWR U$$3276/X sky130_fd_sc_hd__xor2_1
XU$$2531 U$$2531/A U$$2533/B VGND VGND VPWR VPWR U$$2531/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$58 _482_/Q _354_/Q VGND VGND VPWR VPWR final_adder.U$$553/B1 final_adder.U$$680/A
+ sky130_fd_sc_hd__ha_1
XU$$2542 _586_/Q U$$2584/A2 _587_/Q U$$2584/B2 VGND VGND VPWR VPWR U$$2543/A sky130_fd_sc_hd__a22o_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$69 _493_/Q _365_/Q VGND VGND VPWR VPWR final_adder.U$$197/B1 final_adder.U$$691/A
+ sky130_fd_sc_hd__ha_1
XU$$3287 _663_/Q VGND VGND VPWR VPWR U$$3287/Y sky130_fd_sc_hd__inv_1
XU$$3298 U$$969/A1 U$$3412/A2 U$$12/A1 U$$3412/B2 VGND VGND VPWR VPWR U$$3299/A sky130_fd_sc_hd__a22o_1
XU$$2553 U$$2553/A U$$2585/B VGND VGND VPWR VPWR U$$2553/X sky130_fd_sc_hd__xor2_1
XU$$2564 U$$96/B1 U$$2584/A2 U$$785/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2565/A sky130_fd_sc_hd__a22o_1
XFILLER_34_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2575 U$$2575/A _653_/Q VGND VGND VPWR VPWR U$$2575/X sky130_fd_sc_hd__xor2_1
XU$$1830 U$$1830/A U$$1872/B VGND VGND VPWR VPWR U$$1830/X sky130_fd_sc_hd__xor2_1
XU$$1841 U$$4170/A1 U$$1903/A2 U$$3624/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1842/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2586 _608_/Q U$$2470/X _609_/Q U$$2471/X VGND VGND VPWR VPWR U$$2587/A sky130_fd_sc_hd__a22o_1
XU$$1852 U$$1852/A U$$1856/B VGND VGND VPWR VPWR U$$1852/X sky130_fd_sc_hd__xor2_1
XU$$2597 U$$2597/A _653_/Q VGND VGND VPWR VPWR U$$2597/X sky130_fd_sc_hd__xor2_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1863 U$$82/A1 U$$1867/A2 U$$632/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1864/A sky130_fd_sc_hd__a22o_1
XU$$1874 U$$1874/A _643_/Q VGND VGND VPWR VPWR U$$1874/X sky130_fd_sc_hd__xor2_1
XU$$1885 U$$926/A1 U$$1897/A2 _601_/Q U$$1897/B2 VGND VGND VPWR VPWR U$$1886/A sky130_fd_sc_hd__a22o_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1896 U$$1896/A _643_/Q VGND VGND VPWR VPWR U$$1896/X sky130_fd_sc_hd__xor2_1
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_97_0 dadda_fa_5_97_0/A dadda_fa_5_97_0/B dadda_fa_5_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/A dadda_fa_6_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$515 final_adder.U$$642/A final_adder.U$$642/B final_adder.U$$515/B1
+ VGND VGND VPWR VPWR final_adder.U$$643/B sky130_fd_sc_hd__a21o_1
XFILLER_96_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater730 _566_/Q VGND VGND VPWR VPWR U$$36/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$537 final_adder.U$$664/A final_adder.U$$664/B final_adder.U$$537/B1
+ VGND VGND VPWR VPWR final_adder.U$$665/B sky130_fd_sc_hd__a21o_1
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater741 _560_/Q VGND VGND VPWR VPWR U$$983/A1 sky130_fd_sc_hd__buf_12
XFILLER_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater752 _556_/Q VGND VGND VPWR VPWR U$$16/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$559 final_adder.U$$686/A final_adder.U$$686/B final_adder.U$$559/B1
+ VGND VGND VPWR VPWR final_adder.U$$687/B sky130_fd_sc_hd__a21o_1
XU$$409 U$$409/A _621_/Q VGND VGND VPWR VPWR U$$409/X sky130_fd_sc_hd__xor2_1
XFILLER_84_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_106_1 U$$3943/X U$$4076/X U$$4209/X VGND VGND VPWR VPWR dadda_fa_4_107_0/CIN
+ dadda_fa_4_106_2/A sky130_fd_sc_hd__fa_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_785__837 VGND VGND VPWR VPWR _785__837/HI U$$4415/B sky130_fd_sc_hd__conb_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_127_0 U$$4383/Y U$$4517/X input159/X VGND VGND VPWR VPWR dadda_fa_6_127_0/COUT
+ dadda_fa_7_127_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_47_3 dadda_fa_3_47_3/A dadda_fa_3_47_3/B dadda_fa_3_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/B dadda_fa_4_47_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_169_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_826__878 VGND VGND VPWR VPWR _826__878/HI U$$4497/B sky130_fd_sc_hd__conb_1
XFILLER_75_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$910 U$$88/A1 U$$910/A2 U$$90/A1 U$$910/B2 VGND VGND VPWR VPWR U$$911/A sky130_fd_sc_hd__a22o_1
XFILLER_75_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$921 U$$921/A U$$923/B VGND VGND VPWR VPWR U$$921/X sky130_fd_sc_hd__xor2_1
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$932 U$$932/A1 U$$826/X U$$934/A1 U$$827/X VGND VGND VPWR VPWR U$$933/A sky130_fd_sc_hd__a22o_1
XU$$943 U$$943/A U$$943/B VGND VGND VPWR VPWR U$$943/X sky130_fd_sc_hd__xor2_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$954 _614_/Q U$$826/X _615_/Q U$$827/X VGND VGND VPWR VPWR U$$955/A sky130_fd_sc_hd__a22o_1
XU$$1104 _552_/Q U$$1100/X U$$969/A1 U$$1101/X VGND VGND VPWR VPWR U$$1105/A sky130_fd_sc_hd__a22o_1
XU$$965 U$$965/A1 U$$999/A2 U$$8/A1 U$$999/B2 VGND VGND VPWR VPWR U$$966/A sky130_fd_sc_hd__a22o_1
XFILLER_188_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$976 U$$976/A U$$998/B VGND VGND VPWR VPWR U$$976/X sky130_fd_sc_hd__xor2_1
XU$$1115 U$$1115/A U$$1189/B VGND VGND VPWR VPWR U$$1115/X sky130_fd_sc_hd__xor2_1
XFILLER_44_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1126 U$$28/B1 U$$1100/X U$$32/A1 U$$1101/X VGND VGND VPWR VPWR U$$1127/A sky130_fd_sc_hd__a22o_1
XU$$987 U$$987/A1 U$$999/A2 U$$28/B1 U$$987/B2 VGND VGND VPWR VPWR U$$988/A sky130_fd_sc_hd__a22o_1
XU$$1137 U$$1137/A U$$1167/B VGND VGND VPWR VPWR U$$1137/X sky130_fd_sc_hd__xor2_1
XU$$998 U$$998/A U$$998/B VGND VGND VPWR VPWR U$$998/X sky130_fd_sc_hd__xor2_1
XU$$1148 U$$50/B1 U$$1200/A2 U$$876/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1149/A sky130_fd_sc_hd__a22o_1
XU$$1159 U$$1159/A U$$1232/A VGND VGND VPWR VPWR U$$1159/X sky130_fd_sc_hd__xor2_1
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_42_2 U$$2751/X U$$2884/X U$$2996/B VGND VGND VPWR VPWR dadda_fa_3_43_1/A
+ dadda_fa_3_42_3/A sky130_fd_sc_hd__fa_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3040 U$$4273/A1 U$$3090/A2 _562_/Q U$$3090/B2 VGND VGND VPWR VPWR U$$3041/A sky130_fd_sc_hd__a22o_1
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR clkbuf_3_4_0_clk/X sky130_fd_sc_hd__clkbuf_2
XU$$3051 U$$3051/A U$$3109/B VGND VGND VPWR VPWR U$$3051/X sky130_fd_sc_hd__xor2_1
XFILLER_35_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_35_1 U$$742/X U$$875/X U$$1008/X VGND VGND VPWR VPWR dadda_fa_3_36_0/CIN
+ dadda_fa_3_35_2/CIN sky130_fd_sc_hd__fa_1
XU$$3062 _572_/Q U$$3146/A2 U$$735/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3063/A sky130_fd_sc_hd__a22o_1
XU$$3073 U$$3073/A U$$3109/B VGND VGND VPWR VPWR U$$3073/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_0 input160/X dadda_fa_5_12_0/B dadda_fa_5_12_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_6_13_0/A dadda_fa_6_12_0/CIN sky130_fd_sc_hd__fa_2
XU$$3084 U$$892/A1 U$$3090/A2 U$$892/B1 U$$3090/B2 VGND VGND VPWR VPWR U$$3085/A sky130_fd_sc_hd__a22o_1
XU$$3095 U$$3095/A U$$3109/B VGND VGND VPWR VPWR U$$3095/X sky130_fd_sc_hd__xor2_1
XU$$2350 U$$2350/A U$$2432/B VGND VGND VPWR VPWR U$$2350/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_0 U$$63/X U$$196/X U$$329/X VGND VGND VPWR VPWR dadda_fa_3_29_1/CIN
+ dadda_fa_3_28_3/A sky130_fd_sc_hd__fa_2
XU$$2361 U$$30/B1 U$$2333/X U$$34/A1 U$$2334/X VGND VGND VPWR VPWR U$$2362/A sky130_fd_sc_hd__a22o_1
XFILLER_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2372 U$$2372/A U$$2436/B VGND VGND VPWR VPWR U$$2372/X sky130_fd_sc_hd__xor2_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2383 U$$4438/A1 U$$2421/A2 U$$4303/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2384/A
+ sky130_fd_sc_hd__a22o_1
XU$$2394 U$$2394/A U$$2432/B VGND VGND VPWR VPWR U$$2394/X sky130_fd_sc_hd__xor2_1
XU$$1660 U$$16/A1 U$$1734/A2 U$$975/B1 U$$1734/B2 VGND VGND VPWR VPWR U$$1661/A sky130_fd_sc_hd__a22o_1
XU$$1671 U$$1671/A U$$1739/B VGND VGND VPWR VPWR U$$1671/X sky130_fd_sc_hd__xor2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1682 U$$38/A1 U$$1734/A2 U$$3191/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1683/A sky130_fd_sc_hd__a22o_1
XU$$1693 U$$1693/A U$$1727/B VGND VGND VPWR VPWR U$$1693/X sky130_fd_sc_hd__xor2_1
XFILLER_187_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_87_4 U$$3240/X U$$3373/X U$$3506/X VGND VGND VPWR VPWR dadda_fa_2_88_4/B
+ dadda_fa_3_87_0/A sky130_fd_sc_hd__fa_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_57_2 dadda_fa_4_57_2/A dadda_fa_4_57_2/B dadda_fa_4_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/CIN dadda_fa_5_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$301 final_adder.U$$300/A final_adder.U$$217/X final_adder.U$$219/X
+ VGND VGND VPWR VPWR final_adder.U$$301/X sky130_fd_sc_hd__a21o_1
XFILLER_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$312 final_adder.U$$312/A final_adder.U$$312/B VGND VGND VPWR VPWR
+ final_adder.U$$348/B sky130_fd_sc_hd__and2_1
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$323 final_adder.U$$322/A final_adder.U$$261/X final_adder.U$$263/X
+ VGND VGND VPWR VPWR final_adder.U$$323/X sky130_fd_sc_hd__a21o_1
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$334 final_adder.U$$334/A final_adder.U$$334/B VGND VGND VPWR VPWR
+ final_adder.U$$358/A sky130_fd_sc_hd__and2_1
XFILLER_183_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$345 final_adder.U$$344/A final_adder.U$$305/X final_adder.U$$307/X
+ VGND VGND VPWR VPWR final_adder.U$$345/X sky130_fd_sc_hd__a21o_1
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$356 final_adder.U$$356/A final_adder.U$$356/B VGND VGND VPWR VPWR
+ final_adder.U$$370/B sky130_fd_sc_hd__and2_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_27_0 dadda_fa_7_27_0/A dadda_fa_7_27_0/B dadda_fa_7_27_0/CIN VGND VGND
+ VPWR VPWR _452_/D _323_/D sky130_fd_sc_hd__fa_2
Xrepeater560 _651_/Q VGND VGND VPWR VPWR U$$2464/B sky130_fd_sc_hd__buf_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$206 U$$206/A U$$242/B VGND VGND VPWR VPWR U$$206/X sky130_fd_sc_hd__xor2_1
Xrepeater571 _643_/Q VGND VGND VPWR VPWR U$$1918/A sky130_fd_sc_hd__buf_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$217 U$$80/A1 U$$141/X U$$82/A1 U$$142/X VGND VGND VPWR VPWR U$$218/A sky130_fd_sc_hd__a22o_1
Xrepeater582 _637_/Q VGND VGND VPWR VPWR U$$1479/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$389 final_adder.U$$364/X final_adder.U$$718/B final_adder.U$$365/X
+ VGND VGND VPWR VPWR final_adder.U$$734/B sky130_fd_sc_hd__a21o_2
XU$$228 U$$228/A U$$274/A VGND VGND VPWR VPWR U$$228/X sky130_fd_sc_hd__xor2_1
Xrepeater593 U$$959/A VGND VGND VPWR VPWR U$$923/B sky130_fd_sc_hd__buf_12
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$239 U$$924/A1 U$$141/X U$$926/A1 U$$142/X VGND VGND VPWR VPWR U$$240/A sky130_fd_sc_hd__a22o_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_52_1 dadda_fa_3_52_1/A dadda_fa_3_52_1/B dadda_fa_3_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/CIN dadda_fa_4_52_2/A sky130_fd_sc_hd__fa_1
XFILLER_121_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_68_1 U$$675/X U$$808/X U$$941/X VGND VGND VPWR VPWR dadda_fa_1_69_6/A
+ dadda_fa_1_68_7/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_45_0 dadda_fa_3_45_0/A dadda_fa_3_45_0/B dadda_fa_3_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/B dadda_fa_4_45_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$740 U$$740/A U$$778/B VGND VGND VPWR VPWR U$$740/X sky130_fd_sc_hd__xor2_1
XU$$751 U$$66/A1 U$$817/A2 U$$68/A1 U$$785/B2 VGND VGND VPWR VPWR U$$752/A sky130_fd_sc_hd__a22o_1
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_667_ _667_/CLK _667_/D VGND VGND VPWR VPWR _667_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$762 U$$762/A U$$778/B VGND VGND VPWR VPWR U$$762/X sky130_fd_sc_hd__xor2_1
XU$$773 U$$88/A1 U$$785/A2 U$$90/A1 U$$785/B2 VGND VGND VPWR VPWR U$$774/A sky130_fd_sc_hd__a22o_1
XU$$784 U$$784/A U$$784/B VGND VGND VPWR VPWR U$$784/X sky130_fd_sc_hd__xor2_1
XU$$795 U$$932/A1 U$$817/A2 U$$934/A1 U$$817/B2 VGND VGND VPWR VPWR U$$796/A sky130_fd_sc_hd__a22o_1
X_598_ _598_/CLK _598_/D VGND VGND VPWR VPWR _598_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_98_5 U$$4326/X U$$4459/X VGND VGND VPWR VPWR dadda_fa_3_99_2/B dadda_fa_4_98_0/A
+ sky130_fd_sc_hd__ha_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_102_0 dadda_fa_7_102_0/A dadda_fa_7_102_0/B dadda_fa_7_102_0/CIN VGND
+ VGND VPWR VPWR _527_/D _398_/D sky130_fd_sc_hd__fa_2
XFILLER_145_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_97_3 U$$3526/X U$$3659/X U$$3792/X VGND VGND VPWR VPWR dadda_fa_3_98_1/B
+ dadda_fa_3_97_3/B sky130_fd_sc_hd__fa_1
XFILLER_132_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_67_1 dadda_fa_5_67_1/A dadda_fa_5_67_1/B dadda_fa_5_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/B dadda_fa_7_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_113_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_59_8 dadda_fa_1_59_8/A dadda_fa_1_59_8/B dadda_fa_1_59_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_3/A dadda_fa_3_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_55_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_106_0 _696__916/HI U$$3012/X U$$3145/X VGND VGND VPWR VPWR dadda_fa_3_107_3/B
+ dadda_fa_3_106_3/CIN sky130_fd_sc_hd__fa_1
XU$$2180 U$$2180/A U$$2192/A VGND VGND VPWR VPWR U$$2180/X sky130_fd_sc_hd__xor2_1
XFILLER_23_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2191 U$$2192/A VGND VGND VPWR VPWR U$$2191/Y sky130_fd_sc_hd__inv_1
XFILLER_50_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1490 _608_/Q U$$1374/X _609_/Q U$$1375/X VGND VGND VPWR VPWR U$$1491/A sky130_fd_sc_hd__a22o_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_85_1 U$$1906/X U$$2039/X U$$2172/X VGND VGND VPWR VPWR dadda_fa_2_86_2/CIN
+ dadda_fa_2_85_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_62_0 dadda_fa_4_62_0/A dadda_fa_4_62_0/B dadda_fa_4_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/A dadda_fa_5_62_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_0 U$$1227/X U$$1360/X U$$1493/X VGND VGND VPWR VPWR dadda_fa_2_79_0/B
+ dadda_fa_2_78_3/B sky130_fd_sc_hd__fa_2
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$120 _544_/Q _416_/Q VGND VGND VPWR VPWR final_adder.U$$615/B1 final_adder.U$$742/A
+ sky130_fd_sc_hd__ha_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$131 final_adder.U$$625/A final_adder.U$$497/B1 final_adder.U$$3/COUT
+ VGND VGND VPWR VPWR final_adder.U$$131/X sky130_fd_sc_hd__a21o_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3809 U$$4494/A1 U$$3703/X U$$4496/A1 U$$3704/X VGND VGND VPWR VPWR U$$3810/A sky130_fd_sc_hd__a22o_1
XFILLER_73_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$142 final_adder.U$$637/A final_adder.U$$636/A VGND VGND VPWR VPWR
+ final_adder.U$$262/A sky130_fd_sc_hd__and2_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$153 final_adder.U$$647/A final_adder.U$$519/B1 final_adder.U$$153/B1
+ VGND VGND VPWR VPWR final_adder.U$$153/X sky130_fd_sc_hd__a21o_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$164 final_adder.U$$659/A final_adder.U$$658/A VGND VGND VPWR VPWR
+ final_adder.U$$274/B sky130_fd_sc_hd__and2_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$175 final_adder.U$$669/A final_adder.U$$541/B1 final_adder.U$$175/B1
+ VGND VGND VPWR VPWR final_adder.U$$175/X sky130_fd_sc_hd__a21o_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$186 final_adder.U$$681/A final_adder.U$$680/A VGND VGND VPWR VPWR
+ final_adder.U$$284/A sky130_fd_sc_hd__and2_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater390 U$$689/X VGND VGND VPWR VPWR U$$817/A2 sky130_fd_sc_hd__buf_12
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_521_ _537_/CLK _521_/D VGND VGND VPWR VPWR _521_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$197 final_adder.U$$691/A final_adder.U$$563/B1 final_adder.U$$197/B1
+ VGND VGND VPWR VPWR final_adder.U$$197/X sky130_fd_sc_hd__a21o_1
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_452_ _452_/CLK _452_/D VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_383_ _518_/CLK _383_/D VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_77_0 dadda_fa_6_77_0/A dadda_fa_6_77_0/B dadda_fa_6_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_78_0/B dadda_fa_7_77_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput160 c[12] VGND VGND VPWR VPWR input160/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput171 c[22] VGND VGND VPWR VPWR input171/X sky130_fd_sc_hd__buf_2
Xinput182 c[32] VGND VGND VPWR VPWR input182/X sky130_fd_sc_hd__clkbuf_2
Xinput193 c[42] VGND VGND VPWR VPWR input193/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$570 U$$22/A1 U$$626/A2 _560_/Q U$$553/X VGND VGND VPWR VPWR U$$571/A sky130_fd_sc_hd__a22o_1
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$581 U$$581/A U$$661/B VGND VGND VPWR VPWR U$$581/X sky130_fd_sc_hd__xor2_1
XU$$592 _570_/Q U$$626/A2 U$$46/A1 U$$553/X VGND VGND VPWR VPWR U$$593/A sky130_fd_sc_hd__a22o_1
XFILLER_189_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_95_0 U$$2591/X U$$2724/X U$$2857/X VGND VGND VPWR VPWR dadda_fa_3_96_0/B
+ dadda_fa_3_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_71_7 dadda_fa_1_71_7/A dadda_fa_1_71_7/B dadda_fa_1_71_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_2/CIN dadda_fa_2_71_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_64_6 dadda_fa_1_64_6/A dadda_fa_1_64_6/B dadda_fa_1_64_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/B dadda_fa_2_64_5/B sky130_fd_sc_hd__fa_1
XFILLER_189_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_57_5 U$$3180/X U$$3313/X U$$3446/X VGND VGND VPWR VPWR dadda_fa_2_58_2/A
+ dadda_fa_2_57_5/A sky130_fd_sc_hd__fa_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_7_94_0 dadda_fa_7_94_0/A dadda_fa_7_94_0/B dadda_fa_7_94_0/CIN VGND VGND
+ VPWR VPWR _519_/D _390_/D sky130_fd_sc_hd__fa_1
XFILLER_155_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4307 _578_/Q U$$4251/X _579_/Q U$$4252/X VGND VGND VPWR VPWR U$$4308/A sky130_fd_sc_hd__a22o_1
XFILLER_93_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4318 U$$4318/A U$$4384/A VGND VGND VPWR VPWR U$$4318/X sky130_fd_sc_hd__xor2_1
XU$$4329 U$$82/A1 U$$4377/A2 U$$632/A1 U$$4377/B2 VGND VGND VPWR VPWR U$$4330/A sky130_fd_sc_hd__a22o_1
XFILLER_58_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3606 U$$4289/B1 U$$3624/A2 U$$4291/B1 U$$3624/B2 VGND VGND VPWR VPWR U$$3607/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3617 U$$3617/A U$$3698/A VGND VGND VPWR VPWR U$$3617/X sky130_fd_sc_hd__xor2_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3628 _581_/Q U$$3668/A2 U$$4178/A1 U$$3668/B2 VGND VGND VPWR VPWR U$$3629/A sky130_fd_sc_hd__a22o_1
XU$$3639 U$$3639/A U$$3699/A VGND VGND VPWR VPWR U$$3639/X sky130_fd_sc_hd__xor2_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2905 _562_/Q U$$2975/A2 _563_/Q U$$2975/B2 VGND VGND VPWR VPWR U$$2906/A sky130_fd_sc_hd__a22o_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2916 U$$2916/A U$$2960/B VGND VGND VPWR VPWR U$$2916/X sky130_fd_sc_hd__xor2_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2927 U$$735/A1 U$$3009/A2 U$$52/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2928/A sky130_fd_sc_hd__a22o_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2938 U$$2938/A U$$2960/B VGND VGND VPWR VPWR U$$2938/X sky130_fd_sc_hd__xor2_1
X_504_ _510_/CLK _504_/D VGND VGND VPWR VPWR _504_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2949 U$$892/B1 U$$2975/A2 U$$4045/B1 U$$2975/B2 VGND VGND VPWR VPWR U$$2950/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_22_2 U$$1115/X U$$1248/X U$$1381/X VGND VGND VPWR VPWR dadda_fa_4_23_1/A
+ dadda_fa_4_22_2/B sky130_fd_sc_hd__fa_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _454_/CLK _435_/D VGND VGND VPWR VPWR _435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_366_ _366_/CLK _366_/D VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_158_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_297_ _452_/CLK _297_/D VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_5 dadda_fa_2_74_5/A dadda_fa_2_74_5/B dadda_fa_2_74_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_2/A dadda_fa_4_74_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_67_4 dadda_fa_2_67_4/A dadda_fa_2_67_4/B dadda_fa_2_67_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/CIN dadda_fa_3_67_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_104_1 dadda_fa_5_104_1/A dadda_fa_5_104_1/B dadda_fa_5_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/B dadda_fa_7_104_0/A sky130_fd_sc_hd__fa_2
XFILLER_161_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_62_3 U$$3589/X U$$3722/X U$$3855/X VGND VGND VPWR VPWR dadda_fa_2_63_1/B
+ dadda_fa_2_62_4/B sky130_fd_sc_hd__fa_2
XFILLER_41_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_55_2 U$$1580/X U$$1713/X U$$1846/X VGND VGND VPWR VPWR dadda_fa_2_56_1/A
+ dadda_fa_2_55_4/A sky130_fd_sc_hd__fa_1
XFILLER_68_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_32_1 dadda_fa_4_32_1/A dadda_fa_4_32_1/B dadda_fa_4_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/B dadda_fa_5_32_1/B sky130_fd_sc_hd__fa_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_48_1 U$$502/X U$$635/X U$$768/X VGND VGND VPWR VPWR dadda_fa_2_49_1/B
+ dadda_fa_2_48_4/A sky130_fd_sc_hd__fa_2
XFILLER_16_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_25_0 dadda_fa_4_25_0/A dadda_fa_4_25_0/B dadda_fa_4_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/A dadda_fa_5_25_1/A sky130_fd_sc_hd__fa_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_220_ _480_/CLK _220_/D VGND VGND VPWR VPWR _220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_77_3 dadda_fa_3_77_3/A dadda_fa_3_77_3/B dadda_fa_3_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/B dadda_fa_4_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4104 U$$4104/A U$$4109/A VGND VGND VPWR VPWR U$$4104/X sky130_fd_sc_hd__xor2_1
XFILLER_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4115 U$$4113/B _675_/Q _676_/Q U$$4110/Y VGND VGND VPWR VPWR U$$4115/X sky130_fd_sc_hd__a22o_4
XU$$4126 _556_/Q U$$4244/A2 _557_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4127/A sky130_fd_sc_hd__a22o_1
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4137 U$$4137/A U$$4197/B VGND VGND VPWR VPWR U$$4137/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_14_0 U$$35/X U$$168/X VGND VGND VPWR VPWR dadda_fa_4_15_2/B dadda_ha_3_14_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4148 _567_/Q U$$4244/A2 U$$4424/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4149/A sky130_fd_sc_hd__a22o_1
XU$$3403 U$$3403/A U$$3403/B VGND VGND VPWR VPWR U$$3403/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3414 _611_/Q U$$3292/X U$$950/A1 U$$3293/X VGND VGND VPWR VPWR U$$3415/A sky130_fd_sc_hd__a22o_1
XU$$4159 U$$4159/A U$$4247/A VGND VGND VPWR VPWR U$$4159/X sky130_fd_sc_hd__xor2_1
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3425 _665_/Q VGND VGND VPWR VPWR U$$3425/Y sky130_fd_sc_hd__inv_1
XU$$3436 U$$3436/A U$$3496/B VGND VGND VPWR VPWR U$$3436/X sky130_fd_sc_hd__xor2_1
XFILLER_19_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2702 U$$2702/A _655_/Q VGND VGND VPWR VPWR U$$2702/X sky130_fd_sc_hd__xor2_1
XU$$3447 U$$22/A1 U$$3525/A2 U$$4271/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3448/A sky130_fd_sc_hd__a22o_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3458 U$$3458/A U$$3496/B VGND VGND VPWR VPWR U$$3458/X sky130_fd_sc_hd__xor2_1
XU$$2713 U$$4494/A1 U$$2607/X U$$4496/A1 U$$2608/X VGND VGND VPWR VPWR U$$2714/A sky130_fd_sc_hd__a22o_1
XU$$2724 U$$2724/A _655_/Q VGND VGND VPWR VPWR U$$2724/X sky130_fd_sc_hd__xor2_1
XU$$3469 U$$4289/B1 U$$3525/A2 U$$4291/B1 U$$3525/B2 VGND VGND VPWR VPWR U$$3470/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2735 U$$4379/A1 U$$2607/X U$$956/A1 U$$2608/X VGND VGND VPWR VPWR U$$2736/A sky130_fd_sc_hd__a22o_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2746 U$$2746/A1 U$$2796/A2 U$$8/A1 U$$2745/X VGND VGND VPWR VPWR U$$2747/A sky130_fd_sc_hd__a22o_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2757 U$$2757/A U$$2797/B VGND VGND VPWR VPWR U$$2757/X sky130_fd_sc_hd__xor2_1
XFILLER_2_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2768 _562_/Q U$$2796/A2 _563_/Q U$$2834/B2 VGND VGND VPWR VPWR U$$2769/A sky130_fd_sc_hd__a22o_1
XFILLER_15_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2779 U$$2779/A U$$2797/B VGND VGND VPWR VPWR U$$2779/X sky130_fd_sc_hd__xor2_2
XFILLER_178_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_418_ _531_/CLK _418_/D VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_349_ _480_/CLK _349_/D VGND VGND VPWR VPWR _349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_72_2 dadda_fa_2_72_2/A dadda_fa_2_72_2/B dadda_fa_2_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/A dadda_fa_3_72_3/A sky130_fd_sc_hd__fa_2
XFILLER_155_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_65_1 dadda_fa_2_65_1/A dadda_fa_2_65_1/B dadda_fa_2_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/CIN dadda_fa_3_65_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$708 final_adder.U$$708/A final_adder.U$$708/B VGND VGND VPWR VPWR
+ _254_/D sky130_fd_sc_hd__xor2_1
XFILLER_97_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$719 final_adder.U$$719/A final_adder.U$$719/B VGND VGND VPWR VPWR
+ _265_/D sky130_fd_sc_hd__xor2_2
Xdadda_fa_5_42_0 dadda_fa_5_42_0/A dadda_fa_5_42_0/B dadda_fa_5_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/A dadda_fa_6_42_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_58_0 dadda_fa_2_58_0/A dadda_fa_2_58_0/B dadda_fa_2_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/B dadda_fa_3_58_2/B sky130_fd_sc_hd__fa_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3970 U$$819/A1 U$$3970/A2 U$$3970/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3971/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3981 U$$4255/A1 U$$4045/A2 U$$969/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$3982/A
+ sky130_fd_sc_hd__a22o_1
XU$$3992 U$$3992/A U$$4044/B VGND VGND VPWR VPWR U$$3992/X sky130_fd_sc_hd__xor2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_737__789 VGND VGND VPWR VPWR _737__789/HI U$$271/B1 sky130_fd_sc_hd__conb_1
XFILLER_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_87_2 dadda_fa_4_87_2/A dadda_fa_4_87_2/B dadda_fa_4_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/CIN dadda_fa_5_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput261 _271_/Q VGND VGND VPWR VPWR o[103] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_57_0 dadda_fa_7_57_0/A dadda_fa_7_57_0/B dadda_fa_7_57_0/CIN VGND VGND
+ VPWR VPWR _482_/D _353_/D sky130_fd_sc_hd__fa_1
Xoutput272 _281_/Q VGND VGND VPWR VPWR o[113] sky130_fd_sc_hd__buf_2
XFILLER_161_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput283 _291_/Q VGND VGND VPWR VPWR o[123] sky130_fd_sc_hd__buf_2
XFILLER_88_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput294 _186_/Q VGND VGND VPWR VPWR o[18] sky130_fd_sc_hd__buf_2
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_60_0 U$$1989/X U$$2122/X U$$2255/X VGND VGND VPWR VPWR dadda_fa_2_61_0/B
+ dadda_fa_2_60_3/B sky130_fd_sc_hd__fa_2
XFILLER_102_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2009 U$$2009/A U$$2023/B VGND VGND VPWR VPWR U$$2009/X sky130_fd_sc_hd__xor2_1
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1308 U$$1308/A U$$1369/A VGND VGND VPWR VPWR U$$1308/X sky130_fd_sc_hd__xor2_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1319 U$$908/A1 U$$1367/A2 U$$88/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1320/A sky130_fd_sc_hd__a22o_1
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_203_ _333_/CLK _203_/D VGND VGND VPWR VPWR _203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_1 dadda_fa_3_82_1/A dadda_fa_3_82_1/B dadda_fa_3_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/CIN dadda_fa_4_82_2/A sky130_fd_sc_hd__fa_1
XFILLER_125_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_75_0 dadda_fa_3_75_0/A dadda_fa_3_75_0/B dadda_fa_3_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/B dadda_fa_4_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_686__906 VGND VGND VPWR VPWR _686__906/HI _686__906/LO sky130_fd_sc_hd__conb_1
XFILLER_151_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3200 U$$3200/A U$$3224/B VGND VGND VPWR VPWR U$$3200/X sky130_fd_sc_hd__xor2_1
XU$$3211 U$$4170/A1 U$$3243/A2 U$$3624/A1 U$$3243/B2 VGND VGND VPWR VPWR U$$3212/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3222 U$$3222/A U$$3244/B VGND VGND VPWR VPWR U$$3222/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_111_1 dadda_fa_4_111_1/A dadda_fa_4_111_1/B dadda_fa_4_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/B dadda_fa_5_111_1/B sky130_fd_sc_hd__fa_1
XFILLER_4_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3233 _589_/Q U$$3155/X _590_/Q U$$3156/X VGND VGND VPWR VPWR U$$3234/A sky130_fd_sc_hd__a22o_1
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$15 _439_/Q _311_/Q VGND VGND VPWR VPWR final_adder.U$$143/B1 final_adder.U$$637/A
+ sky130_fd_sc_hd__ha_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3244 U$$3244/A U$$3244/B VGND VGND VPWR VPWR U$$3244/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$26 _450_/Q _322_/Q VGND VGND VPWR VPWR final_adder.U$$521/B1 final_adder.U$$648/A
+ sky130_fd_sc_hd__ha_1
XU$$2510 U$$4289/B1 U$$2534/A2 U$$4291/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2511/A
+ sky130_fd_sc_hd__a22o_1
XU$$3255 _600_/Q U$$3155/X U$$928/A1 U$$3156/X VGND VGND VPWR VPWR U$$3256/A sky130_fd_sc_hd__a22o_1
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$37 _461_/Q _333_/Q VGND VGND VPWR VPWR final_adder.U$$165/B1 final_adder.U$$659/A
+ sky130_fd_sc_hd__ha_1
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_104_0 dadda_fa_4_104_0/A dadda_fa_4_104_0/B dadda_fa_4_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/A dadda_fa_5_104_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_37_5 dadda_fa_2_37_5/A dadda_fa_2_37_5/B dadda_fa_2_37_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_38_2/A dadda_fa_4_37_0/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$48 _472_/Q _344_/Q VGND VGND VPWR VPWR final_adder.U$$543/B1 final_adder.U$$670/A
+ sky130_fd_sc_hd__ha_1
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3266 U$$3266/A U$$3270/B VGND VGND VPWR VPWR U$$3266/X sky130_fd_sc_hd__xor2_1
XU$$2521 U$$2521/A U$$2585/B VGND VGND VPWR VPWR U$$2521/X sky130_fd_sc_hd__xor2_1
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3277 _611_/Q U$$3155/X U$$950/A1 U$$3156/X VGND VGND VPWR VPWR U$$3278/A sky130_fd_sc_hd__a22o_1
XU$$2532 U$$66/A1 U$$2574/A2 U$$68/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2533/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$59 _483_/Q _355_/Q VGND VGND VPWR VPWR final_adder.U$$187/B1 final_adder.U$$681/A
+ sky130_fd_sc_hd__ha_1
XU$$2543 U$$2543/A U$$2585/B VGND VGND VPWR VPWR U$$2543/X sky130_fd_sc_hd__xor2_1
XU$$3288 _663_/Q VGND VGND VPWR VPWR U$$3288/Y sky130_fd_sc_hd__inv_1
XFILLER_185_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2554 U$$4335/A1 U$$2470/X _593_/Q U$$2471/X VGND VGND VPWR VPWR U$$2555/A sky130_fd_sc_hd__a22o_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3299 U$$3299/A U$$3413/B VGND VGND VPWR VPWR U$$3299/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1820 U$$1820/A U$$1872/B VGND VGND VPWR VPWR U$$1820/X sky130_fd_sc_hd__xor2_1
XU$$2565 U$$2565/A U$$2585/B VGND VGND VPWR VPWR U$$2565/X sky130_fd_sc_hd__xor2_1
XU$$1831 U$$50/A1 U$$1897/A2 U$$50/B1 U$$1897/B2 VGND VGND VPWR VPWR U$$1832/A sky130_fd_sc_hd__a22o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2576 U$$4494/A1 U$$2584/A2 U$$4496/A1 U$$2584/B2 VGND VGND VPWR VPWR U$$2577/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1842 U$$1842/A U$$1856/B VGND VGND VPWR VPWR U$$1842/X sky130_fd_sc_hd__xor2_1
XU$$2587 U$$2587/A U$$2603/A VGND VGND VPWR VPWR U$$2587/X sky130_fd_sc_hd__xor2_1
XU$$1853 _584_/Q U$$1903/A2 U$$4045/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1854/A sky130_fd_sc_hd__a22o_1
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2598 _614_/Q U$$2470/X U$$956/A1 U$$2471/X VGND VGND VPWR VPWR U$$2599/A sky130_fd_sc_hd__a22o_1
XU$$1864 U$$1864/A U$$1918/A VGND VGND VPWR VPWR U$$1864/X sky130_fd_sc_hd__xor2_1
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1875 U$$94/A1 U$$1785/X U$$94/B1 U$$1786/X VGND VGND VPWR VPWR U$$1876/A sky130_fd_sc_hd__a22o_1
XU$$1886 U$$1886/A U$$1904/B VGND VGND VPWR VPWR U$$1886/X sky130_fd_sc_hd__xor2_1
XFILLER_187_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1897 U$$938/A1 U$$1897/A2 _607_/Q U$$1897/B2 VGND VGND VPWR VPWR U$$1898/A sky130_fd_sc_hd__a22o_1
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_97_1 dadda_fa_5_97_1/A dadda_fa_5_97_1/B dadda_fa_5_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/B dadda_fa_7_97_0/A sky130_fd_sc_hd__fa_2
XFILLER_147_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$505 final_adder.U$$632/A final_adder.U$$632/B final_adder.U$$505/B1
+ VGND VGND VPWR VPWR final_adder.U$$633/B sky130_fd_sc_hd__a21o_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater720 U$$4291/A1 VGND VGND VPWR VPWR U$$4289/B1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$527 final_adder.U$$654/A final_adder.U$$654/B final_adder.U$$527/B1
+ VGND VGND VPWR VPWR final_adder.U$$655/B sky130_fd_sc_hd__a21o_1
Xrepeater731 _565_/Q VGND VGND VPWR VPWR U$$3457/B1 sky130_fd_sc_hd__buf_12
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater742 _560_/Q VGND VGND VPWR VPWR U$$4271/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$549 final_adder.U$$676/A final_adder.U$$676/B final_adder.U$$549/B1
+ VGND VGND VPWR VPWR final_adder.U$$677/B sky130_fd_sc_hd__a21o_1
XFILLER_38_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater753 _555_/Q VGND VGND VPWR VPWR U$$12/B1 sky130_fd_sc_hd__buf_12
XFILLER_72_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4490 U$$654/A1 U$$4388/X U$$4492/A1 U$$4389/X VGND VGND VPWR VPWR U$$4491/A sky130_fd_sc_hd__a22o_2
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_92_0 dadda_fa_4_92_0/A dadda_fa_4_92_0/B dadda_fa_4_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/A dadda_fa_5_92_1/A sky130_fd_sc_hd__fa_1
XFILLER_109_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_106_2 U$$4342/X U$$4475/X input136/X VGND VGND VPWR VPWR dadda_fa_4_107_1/A
+ dadda_fa_4_106_2/B sky130_fd_sc_hd__fa_2
XFILLER_107_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$900 U$$76/B1 U$$910/A2 U$$902/A1 U$$910/B2 VGND VGND VPWR VPWR U$$901/A sky130_fd_sc_hd__a22o_1
XU$$911 U$$911/A U$$923/B VGND VGND VPWR VPWR U$$911/X sky130_fd_sc_hd__xor2_1
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$922 U$$98/B1 U$$928/A2 U$$924/A1 U$$928/B2 VGND VGND VPWR VPWR U$$923/A sky130_fd_sc_hd__a22o_1
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$933 U$$933/A U$$959/A VGND VGND VPWR VPWR U$$933/X sky130_fd_sc_hd__xor2_1
XU$$944 U$$944/A1 U$$826/X U$$946/A1 U$$827/X VGND VGND VPWR VPWR U$$945/A sky130_fd_sc_hd__a22o_1
XFILLER_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$955 U$$955/A _629_/Q VGND VGND VPWR VPWR U$$955/X sky130_fd_sc_hd__xor2_1
XU$$1105 U$$1105/A U$$1189/B VGND VGND VPWR VPWR U$$1105/X sky130_fd_sc_hd__xor2_1
XFILLER_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$966 U$$966/A U$$992/B VGND VGND VPWR VPWR U$$966/X sky130_fd_sc_hd__xor2_1
XFILLER_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1116 U$$20/A1 U$$1200/A2 _559_/Q U$$1200/B2 VGND VGND VPWR VPWR U$$1117/A sky130_fd_sc_hd__a22o_1
XU$$977 U$$18/A1 U$$999/A2 U$$20/A1 U$$999/B2 VGND VGND VPWR VPWR U$$978/A sky130_fd_sc_hd__a22o_1
XU$$1127 U$$1127/A U$$1189/B VGND VGND VPWR VPWR U$$1127/X sky130_fd_sc_hd__xor2_1
XU$$988 U$$988/A U$$992/B VGND VGND VPWR VPWR U$$988/X sky130_fd_sc_hd__xor2_1
XU$$999 U$$40/A1 U$$999/A2 _569_/Q U$$999/B2 VGND VGND VPWR VPWR U$$999/X sky130_fd_sc_hd__a22o_1
XU$$1138 U$$3876/B1 U$$1200/A2 U$$4291/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1139/A
+ sky130_fd_sc_hd__a22o_1
XU$$1149 U$$1149/A U$$1167/B VGND VGND VPWR VPWR U$$1149/X sky130_fd_sc_hd__xor2_1
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_29_3 U$$1262/X U$$1395/X VGND VGND VPWR VPWR dadda_fa_3_30_2/B dadda_fa_4_29_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_42_3 input193/X dadda_fa_2_42_3/B dadda_fa_2_42_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_43_1/B dadda_fa_3_42_3/B sky130_fd_sc_hd__fa_2
XU$$3030 U$$16/A1 U$$3146/A2 U$$975/B1 U$$3146/B2 VGND VGND VPWR VPWR U$$3031/A sky130_fd_sc_hd__a22o_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3041 U$$3041/A U$$3085/B VGND VGND VPWR VPWR U$$3041/X sky130_fd_sc_hd__xor2_1
XFILLER_47_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3052 U$$4285/A1 U$$3090/A2 U$$4424/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3053/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3063 U$$3063/A U$$3129/B VGND VGND VPWR VPWR U$$3063/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_2 U$$1141/X U$$1274/X U$$1407/X VGND VGND VPWR VPWR dadda_fa_3_36_1/A
+ dadda_fa_3_35_3/A sky130_fd_sc_hd__fa_1
XU$$3074 U$$4170/A1 U$$3090/A2 U$$3624/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3075/A
+ sky130_fd_sc_hd__a22o_1
XU$$2340 U$$2340/A U$$2436/B VGND VGND VPWR VPWR U$$2340/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_1 dadda_fa_5_12_1/A dadda_fa_5_12_1/B dadda_ha_4_12_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_13_0/B dadda_fa_7_12_0/A sky130_fd_sc_hd__fa_1
XU$$3085 U$$3085/A U$$3085/B VGND VGND VPWR VPWR U$$3085/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_1 U$$462/X U$$595/X U$$728/X VGND VGND VPWR VPWR dadda_fa_3_29_2/A
+ dadda_fa_3_28_3/B sky130_fd_sc_hd__fa_1
XU$$2351 U$$979/B1 U$$2421/A2 U$$983/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2352/A sky130_fd_sc_hd__a22o_1
XU$$3096 U$$902/B1 U$$3146/A2 _590_/Q U$$3146/B2 VGND VGND VPWR VPWR U$$3097/A sky130_fd_sc_hd__a22o_1
XU$$2362 U$$2362/A U$$2432/B VGND VGND VPWR VPWR U$$2362/X sky130_fd_sc_hd__xor2_1
XU$$2373 U$$4289/B1 U$$2421/A2 U$$4291/B1 U$$2421/B2 VGND VGND VPWR VPWR U$$2374/A
+ sky130_fd_sc_hd__a22o_1
XU$$2384 U$$2384/A U$$2436/B VGND VGND VPWR VPWR U$$2384/X sky130_fd_sc_hd__xor2_1
XU$$1650 U$$1650/A1 U$$1734/A2 U$$8/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1651/A sky130_fd_sc_hd__a22o_1
XU$$2395 U$$66/A1 U$$2333/X _582_/Q U$$2334/X VGND VGND VPWR VPWR U$$2396/A sky130_fd_sc_hd__a22o_1
XU$$1661 U$$1661/A U$$1781/A VGND VGND VPWR VPWR U$$1661/X sky130_fd_sc_hd__xor2_1
XU$$1672 U$$987/A1 U$$1726/A2 U$$30/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1673/A sky130_fd_sc_hd__a22o_1
XU$$1683 U$$1683/A U$$1727/B VGND VGND VPWR VPWR U$$1683/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1694 U$$50/A1 U$$1726/A2 U$$2790/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1695/A sky130_fd_sc_hd__a22o_1
XFILLER_188_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$302 final_adder.U$$302/A final_adder.U$$302/B VGND VGND VPWR VPWR
+ final_adder.U$$342/A sky130_fd_sc_hd__and2_1
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$313 final_adder.U$$312/A final_adder.U$$241/X final_adder.U$$243/X
+ VGND VGND VPWR VPWR final_adder.U$$313/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$324 final_adder.U$$324/A final_adder.U$$324/B VGND VGND VPWR VPWR
+ final_adder.U$$354/B sky130_fd_sc_hd__and2_1
XFILLER_85_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$335 final_adder.U$$334/A final_adder.U$$285/X final_adder.U$$287/X
+ VGND VGND VPWR VPWR final_adder.U$$335/X sky130_fd_sc_hd__a21o_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$346 final_adder.U$$346/A final_adder.U$$346/B VGND VGND VPWR VPWR
+ final_adder.U$$364/A sky130_fd_sc_hd__and2_1
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater550 _657_/Q VGND VGND VPWR VPWR U$$2871/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$357 final_adder.U$$356/A final_adder.U$$329/X final_adder.U$$331/X
+ VGND VGND VPWR VPWR final_adder.U$$357/X sky130_fd_sc_hd__a21o_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater561 U$$2289/B VGND VGND VPWR VPWR U$$2257/B sky130_fd_sc_hd__buf_12
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$207 U$$68/B1 U$$141/X U$$72/A1 U$$142/X VGND VGND VPWR VPWR U$$208/A sky130_fd_sc_hd__a22o_1
Xrepeater572 U$$1872/B VGND VGND VPWR VPWR U$$1856/B sky130_fd_sc_hd__buf_12
XU$$218 U$$218/A U$$242/B VGND VGND VPWR VPWR U$$218/X sky130_fd_sc_hd__xor2_1
Xrepeater583 _637_/Q VGND VGND VPWR VPWR U$$1505/B sky130_fd_sc_hd__buf_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$229 U$$92/A1 U$$141/X U$$92/B1 U$$142/X VGND VGND VPWR VPWR U$$230/A sky130_fd_sc_hd__a22o_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater594 U$$943/B VGND VGND VPWR VPWR U$$903/B sky130_fd_sc_hd__buf_12
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_752__804 VGND VGND VPWR VPWR _752__804/HI U$$3568/A1 sky130_fd_sc_hd__conb_1
XFILLER_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_111_0 U$$3287/Y U$$3421/X U$$3554/X VGND VGND VPWR VPWR dadda_fa_4_112_1/A
+ dadda_fa_4_111_2/A sky130_fd_sc_hd__fa_1
XFILLER_5_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_52_2 dadda_fa_3_52_2/A dadda_fa_3_52_2/B dadda_fa_3_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/A dadda_fa_4_52_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_2 U$$1074/X U$$1207/X U$$1340/X VGND VGND VPWR VPWR dadda_fa_1_69_6/B
+ dadda_fa_1_68_8/A sky130_fd_sc_hd__fa_1
XFILLER_121_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_45_1 dadda_fa_3_45_1/A dadda_fa_3_45_1/B dadda_fa_3_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/CIN dadda_fa_4_45_2/A sky130_fd_sc_hd__fa_2
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_22_0 dadda_fa_6_22_0/A dadda_fa_6_22_0/B dadda_fa_6_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_23_0/B dadda_fa_7_22_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_21_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_38_0 dadda_fa_3_38_0/A dadda_fa_3_38_0/B dadda_fa_3_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/B dadda_fa_4_38_1/CIN sky130_fd_sc_hd__fa_1
XU$$730 U$$730/A U$$784/B VGND VGND VPWR VPWR U$$730/X sky130_fd_sc_hd__xor2_1
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_666_ _669_/CLK _666_/D VGND VGND VPWR VPWR _666_/Q sky130_fd_sc_hd__dfxtp_1
XU$$741 U$$878/A1 U$$785/A2 U$$58/A1 U$$785/B2 VGND VGND VPWR VPWR U$$742/A sky130_fd_sc_hd__a22o_1
XFILLER_189_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$752 U$$752/A U$$784/B VGND VGND VPWR VPWR U$$752/X sky130_fd_sc_hd__xor2_1
XU$$763 U$$76/B1 U$$785/A2 U$$902/A1 U$$785/B2 VGND VGND VPWR VPWR U$$764/A sky130_fd_sc_hd__a22o_1
XU$$774 U$$774/A U$$778/B VGND VGND VPWR VPWR U$$774/X sky130_fd_sc_hd__xor2_1
XFILLER_17_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_597_ _597_/CLK _597_/D VGND VGND VPWR VPWR _597_/Q sky130_fd_sc_hd__dfxtp_4
XU$$785 U$$785/A1 U$$785/A2 U$$924/A1 U$$785/B2 VGND VGND VPWR VPWR U$$786/A sky130_fd_sc_hd__a22o_1
XU$$796 U$$796/A U$$822/A VGND VGND VPWR VPWR U$$796/X sky130_fd_sc_hd__xor2_1
XFILLER_188_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_97_4 U$$3925/X U$$4058/X U$$4191/X VGND VGND VPWR VPWR dadda_fa_3_98_1/CIN
+ dadda_fa_3_97_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_40_0 U$$1550/X U$$1683/X U$$1816/X VGND VGND VPWR VPWR dadda_fa_3_41_0/B
+ dadda_fa_3_40_2/B sky130_fd_sc_hd__fa_2
XFILLER_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2170 U$$2170/A U$$2192/A VGND VGND VPWR VPWR U$$2170/X sky130_fd_sc_hd__xor2_1
XU$$2181 U$$4510/A1 U$$2189/A2 _612_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2182/A sky130_fd_sc_hd__a22o_1
XU$$2192 U$$2192/A VGND VGND VPWR VPWR U$$2192/Y sky130_fd_sc_hd__inv_1
XU$$1480 U$$932/A1 U$$1374/X U$$934/A1 U$$1375/X VGND VGND VPWR VPWR U$$1481/A sky130_fd_sc_hd__a22o_1
XU$$1491 U$$1491/A U$$1505/B VGND VGND VPWR VPWR U$$1491/X sky130_fd_sc_hd__xor2_1
XFILLER_50_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_85_2 U$$2305/X U$$2438/X U$$2571/X VGND VGND VPWR VPWR dadda_fa_2_86_3/A
+ dadda_fa_2_85_5/A sky130_fd_sc_hd__fa_1
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_62_1 dadda_fa_4_62_1/A dadda_fa_4_62_1/B dadda_fa_4_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/B dadda_fa_5_62_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_1 U$$1626/X U$$1759/X U$$1892/X VGND VGND VPWR VPWR dadda_fa_2_79_0/CIN
+ dadda_fa_2_78_3/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_4_55_0 dadda_fa_4_55_0/A dadda_fa_4_55_0/B dadda_fa_4_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/A dadda_fa_5_55_1/A sky130_fd_sc_hd__fa_1
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$110 _534_/Q _406_/Q VGND VGND VPWR VPWR final_adder.U$$605/B1 final_adder.U$$732/A
+ sky130_fd_sc_hd__ha_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$121 _545_/Q _417_/Q VGND VGND VPWR VPWR final_adder.U$$249/B1 final_adder.U$$743/A
+ sky130_fd_sc_hd__ha_1
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$132 final_adder.U$$627/A final_adder.U$$626/A VGND VGND VPWR VPWR
+ final_adder.U$$258/B sky130_fd_sc_hd__and2_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$143 final_adder.U$$637/A final_adder.U$$509/B1 final_adder.U$$143/B1
+ VGND VGND VPWR VPWR final_adder.U$$143/X sky130_fd_sc_hd__a21o_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$154 final_adder.U$$649/A final_adder.U$$648/A VGND VGND VPWR VPWR
+ final_adder.U$$268/A sky130_fd_sc_hd__and2_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$165 final_adder.U$$659/A final_adder.U$$531/B1 final_adder.U$$165/B1
+ VGND VGND VPWR VPWR final_adder.U$$165/X sky130_fd_sc_hd__a21o_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$176 final_adder.U$$671/A final_adder.U$$670/A VGND VGND VPWR VPWR
+ final_adder.U$$280/B sky130_fd_sc_hd__and2_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_520_ _583_/CLK _520_/D VGND VGND VPWR VPWR _520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$187 final_adder.U$$681/A final_adder.U$$553/B1 final_adder.U$$187/B1
+ VGND VGND VPWR VPWR final_adder.U$$187/X sky130_fd_sc_hd__a21o_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater391 U$$626/A2 VGND VGND VPWR VPWR U$$682/A2 sky130_fd_sc_hd__buf_12
XFILLER_79_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$198 final_adder.U$$693/A final_adder.U$$692/A VGND VGND VPWR VPWR
+ final_adder.U$$290/A sky130_fd_sc_hd__and2_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_451_ _458_/CLK _451_/D VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_382_ _387_/CLK _382_/D VGND VGND VPWR VPWR _382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR _369_/CLK sky130_fd_sc_hd__clkbuf_2
Xdadda_ha_0_74_2 U$$1485/X U$$1618/X VGND VGND VPWR VPWR dadda_fa_1_75_8/B dadda_fa_2_74_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_73_0 U$$684/Y U$$818/X U$$951/X VGND VGND VPWR VPWR dadda_fa_1_74_7/B
+ dadda_fa_1_73_8/B sky130_fd_sc_hd__fa_2
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput150 c[119] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput161 c[13] VGND VGND VPWR VPWR input161/X sky130_fd_sc_hd__clkbuf_2
Xinput172 c[23] VGND VGND VPWR VPWR input172/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput183 c[33] VGND VGND VPWR VPWR input183/X sky130_fd_sc_hd__clkbuf_1
Xinput194 c[43] VGND VGND VPWR VPWR input194/X sky130_fd_sc_hd__buf_2
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$560 U$$971/A1 U$$626/A2 U$$12/B1 U$$553/X VGND VGND VPWR VPWR U$$561/A sky130_fd_sc_hd__a22o_1
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_649_ _649_/CLK _649_/D VGND VGND VPWR VPWR _649_/Q sky130_fd_sc_hd__dfxtp_4
XU$$571 U$$571/A U$$623/B VGND VGND VPWR VPWR U$$571/X sky130_fd_sc_hd__xor2_1
XFILLER_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$582 U$$34/A1 U$$626/A2 U$$36/A1 U$$553/X VGND VGND VPWR VPWR U$$583/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$593 U$$593/A U$$623/B VGND VGND VPWR VPWR U$$593/X sky130_fd_sc_hd__xor2_2
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_95_1 U$$2990/X U$$3123/X U$$3256/X VGND VGND VPWR VPWR dadda_fa_3_96_0/CIN
+ dadda_fa_3_95_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_72_0 dadda_fa_5_72_0/A dadda_fa_5_72_0/B dadda_fa_5_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/A dadda_fa_6_72_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_132_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_88_0 U$$3508/X U$$3641/X U$$3774/X VGND VGND VPWR VPWR dadda_fa_3_89_0/B
+ dadda_fa_3_88_2/B sky130_fd_sc_hd__fa_2
XFILLER_114_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_8 dadda_fa_1_71_8/A dadda_fa_1_71_8/B dadda_fa_1_71_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_3/A dadda_fa_3_71_0/A sky130_fd_sc_hd__fa_2
XFILLER_87_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_64_7 dadda_fa_1_64_7/A dadda_fa_1_64_7/B dadda_fa_1_64_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/CIN dadda_fa_2_64_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_57_6 U$$3579/X U$$3712/X U$$3845/X VGND VGND VPWR VPWR dadda_fa_2_58_2/B
+ dadda_fa_2_57_5/B sky130_fd_sc_hd__fa_2
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_9_0 dadda_fa_7_9_0/A dadda_fa_7_9_0/B dadda_fa_7_9_0/CIN VGND VGND VPWR
+ VPWR _434_/D _305_/D sky130_fd_sc_hd__fa_2
XFILLER_39_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_87_0 dadda_fa_7_87_0/A dadda_fa_7_87_0/B dadda_fa_7_87_0/CIN VGND VGND
+ VPWR VPWR _512_/D _383_/D sky130_fd_sc_hd__fa_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_90_0 _690__910/HI U$$1916/X U$$2049/X VGND VGND VPWR VPWR dadda_fa_2_91_4/A
+ dadda_fa_2_90_5/A sky130_fd_sc_hd__fa_2
XFILLER_117_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4308 U$$4308/A U$$4332/B VGND VGND VPWR VPWR U$$4308/X sky130_fd_sc_hd__xor2_1
XU$$4319 _584_/Q U$$4251/X _585_/Q U$$4252/X VGND VGND VPWR VPWR U$$4320/A sky130_fd_sc_hd__a22o_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3607 U$$3607/A U$$3625/B VGND VGND VPWR VPWR U$$3607/X sky130_fd_sc_hd__xor2_1
XU$$3618 U$$4303/A1 U$$3668/A2 _577_/Q U$$3668/B2 VGND VGND VPWR VPWR U$$3619/A sky130_fd_sc_hd__a22o_1
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3629 U$$3629/A U$$3699/A VGND VGND VPWR VPWR U$$3629/X sky130_fd_sc_hd__xor2_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_102_0 dadda_fa_6_102_0/A dadda_fa_6_102_0/B dadda_fa_6_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_103_0/B dadda_fa_7_102_0/CIN sky130_fd_sc_hd__fa_2
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2906 U$$2906/A U$$2960/B VGND VGND VPWR VPWR U$$2906/X sky130_fd_sc_hd__xor2_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2917 U$$4424/A1 U$$2975/A2 U$$4289/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2918/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2928 U$$2928/A U$$2996/B VGND VGND VPWR VPWR U$$2928/X sky130_fd_sc_hd__xor2_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ _503_/CLK _503_/D VGND VGND VPWR VPWR _503_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2939 U$$3624/A1 U$$2975/A2 U$$3900/A1 U$$2975/B2 VGND VGND VPWR VPWR U$$2940/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_22_3 U$$1514/X U$$1614/B input171/X VGND VGND VPWR VPWR dadda_fa_4_23_1/B
+ dadda_fa_4_22_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ _465_/CLK _434_/D VGND VGND VPWR VPWR _434_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_758__810 VGND VGND VPWR VPWR _758__810/HI U$$3979/A1 sky130_fd_sc_hd__conb_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_365_ _366_/CLK _365_/D VGND VGND VPWR VPWR _365_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_296_ _461_/CLK _296_/D VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_67_5 dadda_fa_2_67_5/A dadda_fa_2_67_5/B dadda_fa_2_67_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_2/A dadda_fa_4_67_0/A sky130_fd_sc_hd__fa_2
XFILLER_7_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$390 U$$938/A1 U$$278/X U$$940/A1 U$$279/X VGND VGND VPWR VPWR U$$391/A sky130_fd_sc_hd__a22o_1
XFILLER_177_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_62_4 U$$3988/X U$$4121/X U$$4254/X VGND VGND VPWR VPWR dadda_fa_2_63_1/CIN
+ dadda_fa_2_62_4/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_1_55_3 U$$1979/X U$$2112/X U$$2245/X VGND VGND VPWR VPWR dadda_fa_2_56_1/B
+ dadda_fa_2_55_4/B sky130_fd_sc_hd__fa_2
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_32_2 dadda_fa_4_32_2/A dadda_fa_4_32_2/B dadda_fa_4_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/CIN dadda_fa_5_32_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_2 U$$901/X U$$1034/X U$$1167/X VGND VGND VPWR VPWR dadda_fa_2_49_1/CIN
+ dadda_fa_2_48_4/B sky130_fd_sc_hd__fa_1
XFILLER_83_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_25_1 dadda_fa_4_25_1/A dadda_fa_4_25_1/B dadda_fa_4_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/B dadda_fa_5_25_1/B sky130_fd_sc_hd__fa_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_18_0 U$$1107/X U$$1240/X U$$1336/B VGND VGND VPWR VPWR dadda_fa_5_19_0/A
+ dadda_fa_5_18_1/A sky130_fd_sc_hd__fa_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4105 U$$4379/A1 U$$4107/A2 U$$819/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4106/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4116 U$$4116/A1 U$$4244/A2 _552_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4117/A sky130_fd_sc_hd__a22o_1
XFILLER_120_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4127 U$$4127/A U$$4246/A VGND VGND VPWR VPWR U$$4127/X sky130_fd_sc_hd__xor2_1
XU$$4138 _562_/Q U$$4244/A2 _563_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4139/A sky130_fd_sc_hd__a22o_1
XU$$4149 U$$4149/A U$$4246/A VGND VGND VPWR VPWR U$$4149/X sky130_fd_sc_hd__xor2_1
XU$$3404 _606_/Q U$$3292/X U$$4502/A1 U$$3293/X VGND VGND VPWR VPWR U$$3405/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3415 U$$3415/A _665_/Q VGND VGND VPWR VPWR U$$3415/X sky130_fd_sc_hd__xor2_1
XU$$3426 _666_/Q VGND VGND VPWR VPWR U$$3428/B sky130_fd_sc_hd__inv_1
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3437 U$$4122/A1 U$$3525/A2 U$$14/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3438/A sky130_fd_sc_hd__a22o_1
XFILLER_92_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3448 U$$3448/A U$$3496/B VGND VGND VPWR VPWR U$$3448/X sky130_fd_sc_hd__xor2_1
XFILLER_92_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2703 U$$4484/A1 U$$2607/X _599_/Q U$$2608/X VGND VGND VPWR VPWR U$$2704/A sky130_fd_sc_hd__a22o_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2714 U$$2714/A _655_/Q VGND VGND VPWR VPWR U$$2714/X sky130_fd_sc_hd__xor2_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3459 U$$34/A1 U$$3429/X _566_/Q U$$3430/X VGND VGND VPWR VPWR U$$3460/A sky130_fd_sc_hd__a22o_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2725 _609_/Q U$$2607/X _610_/Q U$$2608/X VGND VGND VPWR VPWR U$$2726/A sky130_fd_sc_hd__a22o_1
XU$$2736 U$$2736/A _655_/Q VGND VGND VPWR VPWR U$$2736/X sky130_fd_sc_hd__xor2_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2747 U$$2747/A U$$2797/B VGND VGND VPWR VPWR U$$2747/X sky130_fd_sc_hd__xor2_2
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_0 U$$47/X U$$180/X U$$313/X VGND VGND VPWR VPWR dadda_fa_4_21_0/B dadda_fa_4_20_1/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2758 U$$4265/A1 U$$2796/A2 U$$979/A1 U$$2826/B2 VGND VGND VPWR VPWR U$$2759/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2769 U$$2769/A U$$2839/B VGND VGND VPWR VPWR U$$2769/X sky130_fd_sc_hd__xor2_1
XFILLER_15_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_417_ _598_/CLK _417_/D VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_348_ _483_/CLK _348_/D VGND VGND VPWR VPWR _348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_279_ _280_/CLK _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_72_3 dadda_fa_2_72_3/A dadda_fa_2_72_3/B dadda_fa_2_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/B dadda_fa_3_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_65_2 dadda_fa_2_65_2/A dadda_fa_2_65_2/B dadda_fa_2_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/A dadda_fa_3_65_3/A sky130_fd_sc_hd__fa_2
XFILLER_64_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$709 final_adder.U$$709/A final_adder.U$$709/B VGND VGND VPWR VPWR
+ _255_/D sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_42_1 dadda_fa_5_42_1/A dadda_fa_5_42_1/B dadda_fa_5_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/B dadda_fa_7_42_0/A sky130_fd_sc_hd__fa_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_58_1 dadda_fa_2_58_1/A dadda_fa_2_58_1/B dadda_fa_2_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/CIN dadda_fa_3_58_2/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_5_35_0 dadda_fa_5_35_0/A dadda_fa_5_35_0/B dadda_fa_5_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/A dadda_fa_6_35_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3960 U$$4508/A1 U$$3970/A2 _611_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3961/A sky130_fd_sc_hd__a22o_1
XU$$3971 U$$3971/A _673_/Q VGND VGND VPWR VPWR U$$3971/X sky130_fd_sc_hd__xor2_1
XU$$3982 U$$3982/A U$$4044/B VGND VGND VPWR VPWR U$$3982/X sky130_fd_sc_hd__xor2_1
XU$$3993 U$$842/A1 U$$4045/A2 _559_/Q U$$4063/B2 VGND VGND VPWR VPWR U$$3994/A sky130_fd_sc_hd__a22o_1
XFILLER_64_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput262 _272_/Q VGND VGND VPWR VPWR o[104] sky130_fd_sc_hd__buf_2
XFILLER_88_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput273 _282_/Q VGND VGND VPWR VPWR o[114] sky130_fd_sc_hd__buf_2
XFILLER_160_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput284 _292_/Q VGND VGND VPWR VPWR o[124] sky130_fd_sc_hd__buf_2
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput295 _187_/Q VGND VGND VPWR VPWR o[19] sky130_fd_sc_hd__buf_2
XFILLER_43_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_60_1 U$$2388/X U$$2521/X U$$2654/X VGND VGND VPWR VPWR dadda_fa_2_61_0/CIN
+ dadda_fa_2_60_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_53_0 U$$379/X U$$512/X U$$645/X VGND VGND VPWR VPWR dadda_fa_2_54_0/B
+ dadda_fa_2_53_3/B sky130_fd_sc_hd__fa_2
XFILLER_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1309 U$$2953/A1 U$$1341/A2 U$$76/B1 U$$1341/B2 VGND VGND VPWR VPWR U$$1310/A sky130_fd_sc_hd__a22o_1
XFILLER_167_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_720__772 VGND VGND VPWR VPWR _720__772/HI U$$1513/A1 sky130_fd_sc_hd__conb_1
XFILLER_169_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_202_ _329_/CLK _202_/D VGND VGND VPWR VPWR _202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_82_2 dadda_fa_3_82_2/A dadda_fa_3_82_2/B dadda_fa_3_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/A dadda_fa_4_82_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_75_1 dadda_fa_3_75_1/A dadda_fa_3_75_1/B dadda_fa_3_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/CIN dadda_fa_4_75_2/A sky130_fd_sc_hd__fa_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_52_0 dadda_fa_6_52_0/A dadda_fa_6_52_0/B dadda_fa_6_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_53_0/B dadda_fa_7_52_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_133_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_68_0 dadda_fa_3_68_0/A dadda_fa_3_68_0/B dadda_fa_3_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/B dadda_fa_4_68_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3201 _573_/Q U$$3241/A2 U$$50/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3202/A sky130_fd_sc_hd__a22o_1
XU$$3212 U$$3212/A U$$3244/B VGND VGND VPWR VPWR U$$3212/X sky130_fd_sc_hd__xor2_1
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_111_2 dadda_fa_4_111_2/A dadda_fa_4_111_2/B dadda_fa_4_111_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/CIN dadda_fa_5_111_1/CIN sky130_fd_sc_hd__fa_2
XU$$3223 U$$72/A1 U$$3241/A2 U$$4045/B1 U$$3253/B2 VGND VGND VPWR VPWR U$$3224/A sky130_fd_sc_hd__a22o_1
XFILLER_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3234 U$$3234/A U$$3270/B VGND VGND VPWR VPWR U$$3234/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$16 _440_/Q _312_/Q VGND VGND VPWR VPWR final_adder.U$$511/B1 final_adder.U$$638/A
+ sky130_fd_sc_hd__ha_1
XFILLER_185_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3245 _595_/Q U$$3155/X _596_/Q U$$3156/X VGND VGND VPWR VPWR U$$3246/A sky130_fd_sc_hd__a22o_1
XU$$2500 U$$3457/B1 U$$2534/A2 U$$4283/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2501/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$27 _451_/Q _323_/Q VGND VGND VPWR VPWR final_adder.U$$155/B1 final_adder.U$$649/A
+ sky130_fd_sc_hd__ha_1
XU$$2511 U$$2511/A U$$2533/B VGND VGND VPWR VPWR U$$2511/X sky130_fd_sc_hd__xor2_1
XU$$3256 U$$3256/A U$$3270/B VGND VGND VPWR VPWR U$$3256/X sky130_fd_sc_hd__xor2_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$38 _462_/Q _334_/Q VGND VGND VPWR VPWR final_adder.U$$533/B1 final_adder.U$$660/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_4_104_1 dadda_fa_4_104_1/A dadda_fa_4_104_1/B dadda_fa_4_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/B dadda_fa_5_104_1/B sky130_fd_sc_hd__fa_1
XU$$3267 U$$4500/A1 U$$3155/X U$$4502/A1 U$$3156/X VGND VGND VPWR VPWR U$$3268/A sky130_fd_sc_hd__a22o_1
XU$$2522 U$$878/A1 U$$2534/A2 U$$880/A1 U$$2534/B2 VGND VGND VPWR VPWR U$$2523/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$49 _473_/Q _345_/Q VGND VGND VPWR VPWR final_adder.U$$177/B1 final_adder.U$$671/A
+ sky130_fd_sc_hd__ha_1
XU$$2533 U$$2533/A U$$2533/B VGND VGND VPWR VPWR U$$2533/X sky130_fd_sc_hd__xor2_1
XU$$3278 U$$3278/A _663_/Q VGND VGND VPWR VPWR U$$3278/X sky130_fd_sc_hd__xor2_1
XU$$2544 _587_/Q U$$2584/A2 _588_/Q U$$2584/B2 VGND VGND VPWR VPWR U$$2545/A sky130_fd_sc_hd__a22o_1
XFILLER_146_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3289 _664_/Q VGND VGND VPWR VPWR U$$3291/B sky130_fd_sc_hd__inv_1
XU$$2555 U$$2555/A U$$2603/A VGND VGND VPWR VPWR U$$2555/X sky130_fd_sc_hd__xor2_1
XU$$1810 U$$1810/A U$$1918/A VGND VGND VPWR VPWR U$$1810/X sky130_fd_sc_hd__xor2_1
XU$$2566 _598_/Q U$$2470/X _599_/Q U$$2471/X VGND VGND VPWR VPWR U$$2567/A sky130_fd_sc_hd__a22o_1
XU$$1821 U$$3191/A1 U$$1897/A2 U$$3876/B1 U$$1897/B2 VGND VGND VPWR VPWR U$$1822/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1832 U$$1832/A U$$1872/B VGND VGND VPWR VPWR U$$1832/X sky130_fd_sc_hd__xor2_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2577 U$$2577/A U$$2603/A VGND VGND VPWR VPWR U$$2577/X sky130_fd_sc_hd__xor2_1
XU$$1843 U$$3624/A1 U$$1903/A2 U$$3900/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1844/A
+ sky130_fd_sc_hd__a22o_1
XU$$2588 U$$4506/A1 U$$2470/X U$$4508/A1 U$$2471/X VGND VGND VPWR VPWR U$$2589/A sky130_fd_sc_hd__a22o_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1854 U$$1854/A U$$1904/B VGND VGND VPWR VPWR U$$1854/X sky130_fd_sc_hd__xor2_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2599 U$$2599/A U$$2603/A VGND VGND VPWR VPWR U$$2599/X sky130_fd_sc_hd__xor2_1
XU$$1865 U$$632/A1 U$$1867/A2 U$$771/A1 U$$1867/B2 VGND VGND VPWR VPWR U$$1866/A sky130_fd_sc_hd__a22o_1
XU$$1876 U$$1876/A U$$1904/B VGND VGND VPWR VPWR U$$1876/X sky130_fd_sc_hd__xor2_1
XFILLER_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1887 U$$654/A1 U$$1785/X U$$930/A1 U$$1786/X VGND VGND VPWR VPWR U$$1888/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_125_0 dadda_fa_7_125_0/A dadda_fa_7_125_0/B dadda_fa_7_125_0/CIN VGND
+ VGND VPWR VPWR _550_/D _421_/D sky130_fd_sc_hd__fa_2
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1898 U$$1898/A U$$1904/B VGND VGND VPWR VPWR U$$1898/X sky130_fd_sc_hd__xor2_1
XFILLER_175_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_70_0 dadda_fa_2_70_0/A dadda_fa_2_70_0/B dadda_fa_2_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/B dadda_fa_3_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater710 U$$50/B1 VGND VGND VPWR VPWR U$$2790/B1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$517 final_adder.U$$644/A final_adder.U$$644/B final_adder.U$$517/B1
+ VGND VGND VPWR VPWR final_adder.U$$645/B sky130_fd_sc_hd__a21o_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater721 _570_/Q VGND VGND VPWR VPWR U$$4291/A1 sky130_fd_sc_hd__buf_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater732 _565_/Q VGND VGND VPWR VPWR U$$34/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$539 final_adder.U$$666/A final_adder.U$$666/B final_adder.U$$539/B1
+ VGND VGND VPWR VPWR final_adder.U$$667/B sky130_fd_sc_hd__a21o_1
Xrepeater743 _559_/Q VGND VGND VPWR VPWR U$$979/B1 sky130_fd_sc_hd__buf_12
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater754 _555_/Q VGND VGND VPWR VPWR U$$14/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4480 U$$94/B1 U$$4388/X U$$98/A1 U$$4389/X VGND VGND VPWR VPWR U$$4481/A sky130_fd_sc_hd__a22o_1
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4491 U$$4491/A U$$4491/B VGND VGND VPWR VPWR U$$4491/X sky130_fd_sc_hd__xor2_4
XFILLER_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3790 U$$3790/A _671_/Q VGND VGND VPWR VPWR U$$3790/X sky130_fd_sc_hd__xor2_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_92_1 dadda_fa_4_92_1/A dadda_fa_4_92_1/B dadda_fa_4_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/B dadda_fa_5_92_1/B sky130_fd_sc_hd__fa_1
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_85_0 dadda_fa_4_85_0/A dadda_fa_4_85_0/B dadda_fa_4_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/A dadda_fa_5_85_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_106_3 dadda_fa_3_106_3/A dadda_fa_3_106_3/B dadda_fa_3_106_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_107_1/B dadda_fa_4_106_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_133_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$901 U$$901/A U$$903/B VGND VGND VPWR VPWR U$$901/X sky130_fd_sc_hd__xor2_1
XU$$912 U$$912/A1 U$$928/A2 U$$914/A1 U$$928/B2 VGND VGND VPWR VPWR U$$913/A sky130_fd_sc_hd__a22o_1
XU$$923 U$$923/A U$$923/B VGND VGND VPWR VPWR U$$923/X sky130_fd_sc_hd__xor2_1
XU$$934 U$$934/A1 U$$826/X U$$936/A1 U$$827/X VGND VGND VPWR VPWR U$$935/A sky130_fd_sc_hd__a22o_1
XU$$945 U$$945/A _629_/Q VGND VGND VPWR VPWR U$$945/X sky130_fd_sc_hd__xor2_1
XFILLER_189_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$956 U$$956/A1 U$$826/X U$$956/B1 U$$827/X VGND VGND VPWR VPWR U$$957/A sky130_fd_sc_hd__a22o_1
XFILLER_141_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$967 _552_/Q U$$963/X U$$969/A1 U$$999/B2 VGND VGND VPWR VPWR U$$968/A sky130_fd_sc_hd__a22o_1
XU$$1106 U$$969/A1 U$$1100/X U$$971/A1 U$$1101/X VGND VGND VPWR VPWR U$$1107/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_82_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _646_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1117 U$$1117/A U$$1189/B VGND VGND VPWR VPWR U$$1117/X sky130_fd_sc_hd__xor2_1
XU$$978 U$$978/A U$$992/B VGND VGND VPWR VPWR U$$978/X sky130_fd_sc_hd__xor2_1
XFILLER_71_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1128 U$$32/A1 U$$1100/X U$$34/A1 U$$1101/X VGND VGND VPWR VPWR U$$1129/A sky130_fd_sc_hd__a22o_1
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$989 U$$28/B1 U$$999/A2 U$$32/A1 U$$999/B2 VGND VGND VPWR VPWR U$$990/A sky130_fd_sc_hd__a22o_1
XU$$1139 U$$1139/A U$$1167/B VGND VGND VPWR VPWR U$$1139/X sky130_fd_sc_hd__xor2_1
XFILLER_44_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3020 U$$3020/A1 U$$3090/A2 U$$4255/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3021/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_42_4 dadda_fa_2_42_4/A dadda_fa_2_42_4/B dadda_fa_2_42_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_1/CIN dadda_fa_3_42_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3031 U$$3031/A U$$3129/B VGND VGND VPWR VPWR U$$3031/X sky130_fd_sc_hd__xor2_1
XFILLER_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3042 U$$28/A1 U$$3146/A2 U$$28/B1 U$$3146/B2 VGND VGND VPWR VPWR U$$3043/A sky130_fd_sc_hd__a22o_1
XFILLER_75_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_35_3 U$$1540/X U$$1673/X U$$1806/X VGND VGND VPWR VPWR dadda_fa_3_36_1/B
+ dadda_fa_3_35_3/B sky130_fd_sc_hd__fa_2
XU$$3053 U$$3053/A U$$3109/B VGND VGND VPWR VPWR U$$3053/X sky130_fd_sc_hd__xor2_1
XFILLER_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3064 U$$735/A1 U$$3146/A2 U$$52/A1 U$$3146/B2 VGND VGND VPWR VPWR U$$3065/A sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3075 U$$3075/A U$$3109/B VGND VGND VPWR VPWR U$$3075/X sky130_fd_sc_hd__xor2_1
XU$$2330 _650_/Q VGND VGND VPWR VPWR U$$2332/B sky130_fd_sc_hd__inv_1
Xclkbuf_leaf_73_clk _560_/CLK VGND VGND VPWR VPWR _576_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3086 U$$892/B1 U$$3146/A2 U$$4045/B1 U$$3146/B2 VGND VGND VPWR VPWR U$$3087/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2341 U$$971/A1 U$$2333/X U$$12/B1 U$$2334/X VGND VGND VPWR VPWR U$$2342/A sky130_fd_sc_hd__a22o_1
XU$$2352 U$$2352/A U$$2432/B VGND VGND VPWR VPWR U$$2352/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_2 U$$861/X U$$994/X U$$1127/X VGND VGND VPWR VPWR dadda_fa_3_29_2/B
+ dadda_fa_3_28_3/CIN sky130_fd_sc_hd__fa_1
XU$$3097 U$$3097/A U$$3109/B VGND VGND VPWR VPWR U$$3097/X sky130_fd_sc_hd__xor2_1
XU$$2363 U$$34/A1 U$$2333/X U$$36/A1 U$$2334/X VGND VGND VPWR VPWR U$$2364/A sky130_fd_sc_hd__a22o_1
XU$$2374 U$$2374/A U$$2436/B VGND VGND VPWR VPWR U$$2374/X sky130_fd_sc_hd__xor2_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2385 U$$4303/A1 U$$2421/A2 U$$4442/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2386/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1640 U$$1640/A _639_/Q VGND VGND VPWR VPWR U$$1640/X sky130_fd_sc_hd__xor2_1
XFILLER_90_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2396 U$$2396/A U$$2464/B VGND VGND VPWR VPWR U$$2396/X sky130_fd_sc_hd__xor2_1
XU$$1651 U$$1651/A U$$1727/B VGND VGND VPWR VPWR U$$1651/X sky130_fd_sc_hd__xor2_1
XU$$1662 U$$975/B1 U$$1734/A2 U$$842/A1 U$$1734/B2 VGND VGND VPWR VPWR U$$1663/A sky130_fd_sc_hd__a22o_1
XU$$1673 U$$1673/A U$$1739/B VGND VGND VPWR VPWR U$$1673/X sky130_fd_sc_hd__xor2_1
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1684 U$$3191/A1 U$$1734/A2 U$$3876/B1 U$$1734/B2 VGND VGND VPWR VPWR U$$1685/A
+ sky130_fd_sc_hd__a22o_1
XU$$1695 U$$1695/A U$$1727/B VGND VGND VPWR VPWR U$$1695/X sky130_fd_sc_hd__xor2_1
XFILLER_33_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$303 final_adder.U$$302/A final_adder.U$$221/X final_adder.U$$223/X
+ VGND VGND VPWR VPWR final_adder.U$$303/X sky130_fd_sc_hd__a21o_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$314 final_adder.U$$314/A final_adder.U$$314/B VGND VGND VPWR VPWR
+ final_adder.U$$348/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$325 final_adder.U$$324/A final_adder.U$$265/X final_adder.U$$267/X
+ VGND VGND VPWR VPWR final_adder.U$$325/X sky130_fd_sc_hd__a21o_1
XFILLER_58_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$336 final_adder.U$$336/A final_adder.U$$336/B VGND VGND VPWR VPWR
+ final_adder.U$$360/B sky130_fd_sc_hd__and2_1
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater540 U$$3270/B VGND VGND VPWR VPWR U$$3244/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$347 final_adder.U$$346/A final_adder.U$$309/X final_adder.U$$311/X
+ VGND VGND VPWR VPWR final_adder.U$$347/X sky130_fd_sc_hd__a21o_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater551 _657_/Q VGND VGND VPWR VPWR U$$2797/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$358 final_adder.U$$358/A final_adder.U$$358/B VGND VGND VPWR VPWR
+ final_adder.U$$370/A sky130_fd_sc_hd__and2_2
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater562 U$$2327/B VGND VGND VPWR VPWR U$$2289/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$369 final_adder.U$$354/X final_adder.U$$638/B final_adder.U$$355/X
+ VGND VGND VPWR VPWR final_adder.U$$654/B sky130_fd_sc_hd__a21o_4
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$208 U$$208/A U$$242/B VGND VGND VPWR VPWR U$$208/X sky130_fd_sc_hd__xor2_1
Xrepeater573 U$$1904/B VGND VGND VPWR VPWR U$$1872/B sky130_fd_sc_hd__buf_12
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$219 U$$82/A1 U$$141/X U$$84/A1 U$$142/X VGND VGND VPWR VPWR U$$220/A sky130_fd_sc_hd__a22o_1
Xrepeater584 U$$1342/B VGND VGND VPWR VPWR U$$1336/B sky130_fd_sc_hd__buf_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater595 U$$959/A VGND VGND VPWR VPWR U$$943/B sky130_fd_sc_hd__buf_12
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_clk clkbuf_3_4_0_clk/X VGND VGND VPWR VPWR _495_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_791__843 VGND VGND VPWR VPWR _791__843/HI U$$4427/B sky130_fd_sc_hd__conb_1
XFILLER_21_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_111_1 U$$3687/X U$$3820/X U$$3953/X VGND VGND VPWR VPWR dadda_fa_4_112_1/B
+ dadda_fa_4_111_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_832__884 VGND VGND VPWR VPWR _832__884/HI U$$4509/B sky130_fd_sc_hd__conb_1
Xdadda_fa_3_104_0 U$$3806/X U$$3939/X U$$4072/X VGND VGND VPWR VPWR dadda_fa_4_105_0/B
+ dadda_fa_4_104_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_52_3 dadda_fa_3_52_3/A dadda_fa_3_52_3/B dadda_fa_3_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/B dadda_fa_4_52_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_3 U$$1473/X U$$1606/X U$$1739/X VGND VGND VPWR VPWR dadda_fa_1_69_6/CIN
+ dadda_fa_1_68_8/B sky130_fd_sc_hd__fa_2
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_45_2 dadda_fa_3_45_2/A dadda_fa_3_45_2/B dadda_fa_3_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/A dadda_fa_4_45_2/B sky130_fd_sc_hd__fa_1
XFILLER_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_38_1 dadda_fa_3_38_1/A dadda_fa_3_38_1/B dadda_fa_3_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/CIN dadda_fa_4_38_2/A sky130_fd_sc_hd__fa_2
X_665_ _669_/CLK _665_/D VGND VGND VPWR VPWR _665_/Q sky130_fd_sc_hd__dfxtp_4
XU$$720 U$$720/A U$$778/B VGND VGND VPWR VPWR U$$720/X sky130_fd_sc_hd__xor2_1
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$731 U$$46/A1 U$$689/X _572_/Q U$$817/B2 VGND VGND VPWR VPWR U$$732/A sky130_fd_sc_hd__a22o_1
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$742 U$$742/A U$$778/B VGND VGND VPWR VPWR U$$742/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_55_clk _536_/CLK VGND VGND VPWR VPWR _598_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_15_0 dadda_fa_6_15_0/A dadda_fa_6_15_0/B dadda_fa_6_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_16_0/B dadda_fa_7_15_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_189_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$753 _582_/Q U$$817/A2 U$$70/A1 U$$785/B2 VGND VGND VPWR VPWR U$$754/A sky130_fd_sc_hd__a22o_1
XU$$764 U$$764/A U$$778/B VGND VGND VPWR VPWR U$$764/X sky130_fd_sc_hd__xor2_1
X_596_ _597_/CLK _596_/D VGND VGND VPWR VPWR _596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$775 U$$912/A1 U$$785/A2 U$$914/A1 U$$785/B2 VGND VGND VPWR VPWR U$$776/A sky130_fd_sc_hd__a22o_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$786 U$$786/A _627_/Q VGND VGND VPWR VPWR U$$786/X sky130_fd_sc_hd__xor2_1
XU$$797 U$$934/A1 U$$689/X U$$799/A1 U$$690/X VGND VGND VPWR VPWR U$$798/A sky130_fd_sc_hd__a22o_1
XFILLER_16_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_3_110_3 U$$4350/X U$$4483/X VGND VGND VPWR VPWR dadda_fa_4_111_1/CIN dadda_ha_3_110_3/SUM
+ sky130_fd_sc_hd__ha_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_97_5 U$$4324/X U$$4457/X input253/X VGND VGND VPWR VPWR dadda_fa_3_98_2/A
+ dadda_fa_4_97_0/A sky130_fd_sc_hd__fa_2
XFILLER_160_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_40_1 U$$1949/X U$$2082/X U$$2215/X VGND VGND VPWR VPWR dadda_fa_3_41_0/CIN
+ dadda_fa_3_40_2/CIN sky130_fd_sc_hd__fa_2
Xclkbuf_leaf_46_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _532_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_33_0 U$$73/X U$$206/X U$$339/X VGND VGND VPWR VPWR dadda_fa_3_34_0/B dadda_fa_3_33_2/B
+ sky130_fd_sc_hd__fa_2
XFILLER_187_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2160 U$$2160/A U$$2192/A VGND VGND VPWR VPWR U$$2160/X sky130_fd_sc_hd__xor2_1
XU$$2171 U$$938/A1 U$$2189/A2 U$$940/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2172/A sky130_fd_sc_hd__a22o_1
XFILLER_179_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2182 U$$2182/A U$$2192/A VGND VGND VPWR VPWR U$$2182/X sky130_fd_sc_hd__xor2_1
XFILLER_168_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2193 _648_/Q VGND VGND VPWR VPWR U$$2195/B sky130_fd_sc_hd__inv_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1470 U$$4484/A1 U$$1374/X _599_/Q U$$1375/X VGND VGND VPWR VPWR U$$1471/A sky130_fd_sc_hd__a22o_1
X_775__827 VGND VGND VPWR VPWR _775__827/HI U$$4395/B sky130_fd_sc_hd__conb_1
XU$$1481 U$$1481/A U$$1505/B VGND VGND VPWR VPWR U$$1481/X sky130_fd_sc_hd__xor2_1
XU$$1492 _609_/Q U$$1374/X _610_/Q U$$1375/X VGND VGND VPWR VPWR U$$1493/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_86_5 U$$3504/X U$$3637/X VGND VGND VPWR VPWR dadda_fa_2_87_4/B dadda_fa_3_86_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_159_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_816__868 VGND VGND VPWR VPWR _816__868/HI U$$4477/B sky130_fd_sc_hd__conb_1
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_85_3 U$$2704/X U$$2837/X U$$2970/X VGND VGND VPWR VPWR dadda_fa_2_86_3/B
+ dadda_fa_2_85_5/B sky130_fd_sc_hd__fa_1
XFILLER_132_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_62_2 dadda_fa_4_62_2/A dadda_fa_4_62_2/B dadda_fa_4_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/CIN dadda_fa_5_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_78_2 U$$2025/X U$$2158/X U$$2291/X VGND VGND VPWR VPWR dadda_fa_2_79_1/A
+ dadda_fa_2_78_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_55_1 dadda_fa_4_55_1/A dadda_fa_4_55_1/B dadda_fa_4_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/B dadda_fa_5_55_1/B sky130_fd_sc_hd__fa_1
XFILLER_98_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$100 _524_/Q _396_/Q VGND VGND VPWR VPWR final_adder.U$$595/B1 final_adder.U$$722/A
+ sky130_fd_sc_hd__ha_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$111 _535_/Q _407_/Q VGND VGND VPWR VPWR final_adder.U$$239/B1 final_adder.U$$733/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_7_32_0 dadda_fa_7_32_0/A dadda_fa_7_32_0/B dadda_fa_7_32_0/CIN VGND VGND
+ VPWR VPWR _457_/D _328_/D sky130_fd_sc_hd__fa_2
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$122 _546_/Q _418_/Q VGND VGND VPWR VPWR final_adder.U$$617/B1 final_adder.U$$744/A
+ sky130_fd_sc_hd__ha_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_0 dadda_fa_4_48_0/A dadda_fa_4_48_0/B dadda_fa_4_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/A dadda_fa_5_48_1/A sky130_fd_sc_hd__fa_1
XFILLER_100_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$133 final_adder.U$$627/A final_adder.U$$499/B1 final_adder.U$$5/COUT
+ VGND VGND VPWR VPWR final_adder.U$$133/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$144 final_adder.U$$639/A final_adder.U$$638/A VGND VGND VPWR VPWR
+ final_adder.U$$264/B sky130_fd_sc_hd__and2_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$155 final_adder.U$$649/A final_adder.U$$521/B1 final_adder.U$$155/B1
+ VGND VGND VPWR VPWR final_adder.U$$155/X sky130_fd_sc_hd__a21o_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$166 final_adder.U$$661/A final_adder.U$$660/A VGND VGND VPWR VPWR
+ final_adder.U$$274/A sky130_fd_sc_hd__and2_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$177 final_adder.U$$671/A final_adder.U$$543/B1 final_adder.U$$177/B1
+ VGND VGND VPWR VPWR final_adder.U$$177/X sky130_fd_sc_hd__a21o_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$188 final_adder.U$$683/A final_adder.U$$682/A VGND VGND VPWR VPWR
+ final_adder.U$$286/B sky130_fd_sc_hd__and2_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater392 U$$552/X VGND VGND VPWR VPWR U$$626/A2 sky130_fd_sc_hd__buf_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$199 final_adder.U$$693/A final_adder.U$$565/B1 final_adder.U$$199/B1
+ VGND VGND VPWR VPWR final_adder.U$$199/X sky130_fd_sc_hd__a21o_1
XFILLER_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _501_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ _462_/CLK _450_/D VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_381_ _510_/CLK _381_/D VGND VGND VPWR VPWR _381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_73_1 U$$1084/X U$$1217/X U$$1350/X VGND VGND VPWR VPWR dadda_fa_1_74_7/CIN
+ dadda_fa_1_73_8/CIN sky130_fd_sc_hd__fa_2
XFILLER_110_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput140 c[10] VGND VGND VPWR VPWR input140/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_50_0 dadda_fa_3_50_0/A dadda_fa_3_50_0/B dadda_fa_3_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/B dadda_fa_4_50_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_76_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_66_0 U$$89/B U$$272/X U$$405/X VGND VGND VPWR VPWR dadda_fa_1_67_5/B dadda_fa_1_66_7/B
+ sky130_fd_sc_hd__fa_1
Xinput151 c[11] VGND VGND VPWR VPWR input151/X sky130_fd_sc_hd__clkbuf_1
Xinput162 c[14] VGND VGND VPWR VPWR input162/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput173 c[24] VGND VGND VPWR VPWR input173/X sky130_fd_sc_hd__buf_2
XFILLER_23_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput184 c[34] VGND VGND VPWR VPWR input184/X sky130_fd_sc_hd__buf_4
XFILLER_36_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput195 c[44] VGND VGND VPWR VPWR input195/X sky130_fd_sc_hd__buf_2
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_clk _369_/CLK VGND VGND VPWR VPWR _490_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$550 _625_/Q VGND VGND VPWR VPWR U$$550/Y sky130_fd_sc_hd__inv_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$561 U$$561/A U$$623/B VGND VGND VPWR VPWR U$$561/X sky130_fd_sc_hd__xor2_1
X_648_ _656_/CLK _648_/D VGND VGND VPWR VPWR _648_/Q sky130_fd_sc_hd__dfxtp_2
XU$$572 U$$983/A1 U$$626/A2 U$$26/A1 U$$553/X VGND VGND VPWR VPWR U$$573/A sky130_fd_sc_hd__a22o_1
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$583 U$$583/A U$$623/B VGND VGND VPWR VPWR U$$583/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$594 U$$46/A1 U$$626/A2 _572_/Q U$$553/X VGND VGND VPWR VPWR U$$595/A sky130_fd_sc_hd__a22o_1
X_579_ _579_/CLK _579_/D VGND VGND VPWR VPWR _579_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_95_2 U$$3389/X U$$3522/X U$$3655/X VGND VGND VPWR VPWR dadda_fa_3_96_1/A
+ dadda_fa_3_95_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_72_1 dadda_fa_5_72_1/A dadda_fa_5_72_1/B dadda_fa_5_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/B dadda_fa_7_72_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_88_1 U$$3907/X U$$4040/X U$$4173/X VGND VGND VPWR VPWR dadda_fa_3_89_0/CIN
+ dadda_fa_3_88_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_65_0 dadda_fa_5_65_0/A dadda_fa_5_65_0/B dadda_fa_5_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/A dadda_fa_6_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_64_8 dadda_fa_1_64_8/A dadda_fa_1_64_8/B dadda_fa_1_64_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_3/A dadda_fa_3_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_57_7 input209/X dadda_fa_1_57_7/B dadda_fa_1_57_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_58_2/CIN dadda_fa_2_57_5/CIN sky130_fd_sc_hd__fa_2
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _448_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_4_0 U$$281/X U$$357/B input201/X VGND VGND VPWR VPWR dadda_fa_7_5_0/B
+ dadda_fa_7_4_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_90_1 U$$2182/X U$$2315/X U$$2448/X VGND VGND VPWR VPWR dadda_fa_2_91_4/B
+ dadda_fa_2_90_5/B sky130_fd_sc_hd__fa_1
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_83_0 U$$1369/Y U$$1503/X U$$1636/X VGND VGND VPWR VPWR dadda_fa_2_84_1/CIN
+ dadda_fa_2_83_4/A sky130_fd_sc_hd__fa_2
XFILLER_89_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4309 U$$4446/A1 U$$4251/X _580_/Q U$$4252/X VGND VGND VPWR VPWR U$$4310/A sky130_fd_sc_hd__a22o_1
XFILLER_58_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3608 U$$4291/B1 U$$3624/A2 U$$4156/B1 U$$3624/B2 VGND VGND VPWR VPWR U$$3609/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3619 U$$3619/A U$$3699/A VGND VGND VPWR VPWR U$$3619/X sky130_fd_sc_hd__xor2_1
XFILLER_73_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2907 _563_/Q U$$2975/A2 _564_/Q U$$2975/B2 VGND VGND VPWR VPWR U$$2908/A sky130_fd_sc_hd__a22o_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2918 U$$2918/A U$$2960/B VGND VGND VPWR VPWR U$$2918/X sky130_fd_sc_hd__xor2_1
XFILLER_34_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ _503_/CLK _502_/D VGND VGND VPWR VPWR _502_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2929 U$$52/A1 U$$3009/A2 U$$54/A1 U$$3009/B2 VGND VGND VPWR VPWR U$$2930/A sky130_fd_sc_hd__a22o_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _465_/CLK _433_/D VGND VGND VPWR VPWR _433_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ _647_/CLK _364_/D VGND VGND VPWR VPWR _364_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_295_ _612_/CLK _295_/D VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_838__890 VGND VGND VPWR VPWR _838__890/HI U$$545/B1 sky130_fd_sc_hd__conb_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_82_0 dadda_fa_6_82_0/A dadda_fa_6_82_0/B dadda_fa_6_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_83_0/B dadda_fa_7_82_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_98_0 input254/X dadda_fa_3_98_0/B dadda_fa_3_98_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_99_0/B dadda_fa_4_98_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_155_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$380 U$$928/A1 U$$278/X U$$930/A1 U$$279/X VGND VGND VPWR VPWR U$$381/A sky130_fd_sc_hd__a22o_1
XFILLER_178_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$391 U$$391/A U$$391/B VGND VGND VPWR VPWR U$$391/X sky130_fd_sc_hd__xor2_1
XFILLER_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk _431_/CLK VGND VGND VPWR VPWR _454_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_5 _679_/Q input215/X dadda_fa_1_62_5/CIN VGND VGND VPWR VPWR dadda_fa_2_63_2/A
+ dadda_fa_2_62_5/A sky130_fd_sc_hd__fa_2
XFILLER_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_4 U$$2378/X U$$2511/X U$$2644/X VGND VGND VPWR VPWR dadda_fa_2_56_1/CIN
+ dadda_fa_2_55_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_48_3 U$$1300/X U$$1433/X U$$1566/X VGND VGND VPWR VPWR dadda_fa_2_49_2/A
+ dadda_fa_2_48_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_4_25_2 dadda_fa_4_25_2/A dadda_fa_4_25_2/B dadda_fa_4_25_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/CIN dadda_fa_5_25_1/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_2_0_clk/X sky130_fd_sc_hd__clkbuf_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_18_1 input166/X dadda_fa_4_18_1/B dadda_fa_4_18_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_19_0/B dadda_fa_5_18_1/B sky130_fd_sc_hd__fa_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4106 U$$4106/A U$$4109/A VGND VGND VPWR VPWR U$$4106/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_21_3 U$$1246/X U$$1379/X VGND VGND VPWR VPWR dadda_fa_4_22_1/B dadda_ha_3_21_3/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4117 U$$4117/A _677_/Q VGND VGND VPWR VPWR U$$4117/X sky130_fd_sc_hd__xor2_1
XU$$4128 _557_/Q U$$4244/A2 _558_/Q U$$4244/B2 VGND VGND VPWR VPWR U$$4129/A sky130_fd_sc_hd__a22o_1
XFILLER_120_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$4139 U$$4139/A _677_/Q VGND VGND VPWR VPWR U$$4139/X sky130_fd_sc_hd__xor2_1
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3405 U$$3405/A _665_/Q VGND VGND VPWR VPWR U$$3405/X sky130_fd_sc_hd__xor2_1
XU$$3416 U$$539/A1 U$$3292/X U$$4514/A1 U$$3293/X VGND VGND VPWR VPWR U$$3417/A sky130_fd_sc_hd__a22o_1
XFILLER_19_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3427 _667_/Q VGND VGND VPWR VPWR U$$3427/Y sky130_fd_sc_hd__inv_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3438 U$$3438/A U$$3496/B VGND VGND VPWR VPWR U$$3438/X sky130_fd_sc_hd__xor2_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3449 U$$4271/A1 U$$3525/A2 U$$4273/A1 U$$3525/B2 VGND VGND VPWR VPWR U$$3450/A
+ sky130_fd_sc_hd__a22o_1
XU$$2704 U$$2704/A _655_/Q VGND VGND VPWR VPWR U$$2704/X sky130_fd_sc_hd__xor2_1
XU$$2715 _604_/Q U$$2607/X _605_/Q U$$2608/X VGND VGND VPWR VPWR U$$2716/A sky130_fd_sc_hd__a22o_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2726 U$$2726/A _655_/Q VGND VGND VPWR VPWR U$$2726/X sky130_fd_sc_hd__xor2_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2737 U$$956/A1 U$$2607/X U$$2737/B1 U$$2608/X VGND VGND VPWR VPWR U$$2738/A sky130_fd_sc_hd__a22o_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_1 U$$446/X U$$579/X U$$712/X VGND VGND VPWR VPWR dadda_fa_4_21_0/CIN
+ dadda_fa_4_20_2/A sky130_fd_sc_hd__fa_2
XU$$2748 U$$8/A1 U$$2796/A2 U$$8/B1 U$$2745/X VGND VGND VPWR VPWR U$$2749/A sky130_fd_sc_hd__a22o_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2759 U$$2759/A U$$2797/B VGND VGND VPWR VPWR U$$2759/X sky130_fd_sc_hd__xor2_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _614_/CLK _416_/D VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_347_ _476_/CLK _347_/D VGND VGND VPWR VPWR _347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_278_ _280_/CLK _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_72_4 dadda_fa_2_72_4/A dadda_fa_2_72_4/B dadda_fa_2_72_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/CIN dadda_fa_3_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_65_3 dadda_fa_2_65_3/A dadda_fa_2_65_3/B dadda_fa_2_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/B dadda_fa_3_65_3/B sky130_fd_sc_hd__fa_1
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_58_2 dadda_fa_2_58_2/A dadda_fa_2_58_2/B dadda_fa_2_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/A dadda_fa_3_58_3/A sky130_fd_sc_hd__fa_2
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_35_1 dadda_fa_5_35_1/A dadda_fa_5_35_1/B dadda_fa_5_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/B dadda_fa_7_35_0/A sky130_fd_sc_hd__fa_1
XFILLER_37_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_28_0 dadda_fa_5_28_0/A dadda_fa_5_28_0/B dadda_fa_5_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/A dadda_fa_6_28_0/CIN sky130_fd_sc_hd__fa_1
XU$$3950 U$$936/A1 U$$3970/A2 U$$4500/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3951/A
+ sky130_fd_sc_hd__a22o_1
XU$$3961 U$$3961/A U$$3969/B VGND VGND VPWR VPWR U$$3961/X sky130_fd_sc_hd__xor2_1
XU$$3972 _673_/Q VGND VGND VPWR VPWR U$$3972/Y sky130_fd_sc_hd__inv_1
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3983 U$$969/A1 U$$4045/A2 U$$12/A1 U$$4063/B2 VGND VGND VPWR VPWR U$$3984/A sky130_fd_sc_hd__a22o_1
XU$$3994 U$$3994/A U$$4044/B VGND VGND VPWR VPWR U$$3994/X sky130_fd_sc_hd__xor2_1
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_102_0 dadda_fa_5_102_0/A dadda_fa_5_102_0/B dadda_fa_5_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/A dadda_fa_6_102_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_134_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput263 _273_/Q VGND VGND VPWR VPWR o[105] sky130_fd_sc_hd__buf_2
Xoutput274 _283_/Q VGND VGND VPWR VPWR o[115] sky130_fd_sc_hd__buf_2
Xoutput285 _293_/Q VGND VGND VPWR VPWR o[125] sky130_fd_sc_hd__buf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput296 _169_/Q VGND VGND VPWR VPWR o[1] sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_60_2 U$$2787/X U$$2920/X U$$3053/X VGND VGND VPWR VPWR dadda_fa_2_61_1/A
+ dadda_fa_2_60_4/A sky130_fd_sc_hd__fa_2
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_53_1 U$$778/X U$$911/X U$$1044/X VGND VGND VPWR VPWR dadda_fa_2_54_0/CIN
+ dadda_fa_2_53_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_30_0 dadda_fa_4_30_0/A dadda_fa_4_30_0/B dadda_fa_4_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/A dadda_fa_5_30_1/A sky130_fd_sc_hd__fa_1
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_46_0 U$$99/X U$$232/X U$$365/X VGND VGND VPWR VPWR dadda_fa_2_47_1/CIN
+ dadda_fa_2_46_4/A sky130_fd_sc_hd__fa_2
XFILLER_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_201_ _456_/CLK _201_/D VGND VGND VPWR VPWR _201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_82_3 dadda_fa_3_82_3/A dadda_fa_3_82_3/B dadda_fa_3_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/B dadda_fa_4_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_75_2 dadda_fa_3_75_2/A dadda_fa_3_75_2/B dadda_fa_3_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/A dadda_fa_4_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_68_1 dadda_fa_3_68_1/A dadda_fa_3_68_1/B dadda_fa_3_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/CIN dadda_fa_4_68_2/A sky130_fd_sc_hd__fa_1
XFILLER_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_45_0 dadda_fa_6_45_0/A dadda_fa_6_45_0/B dadda_fa_6_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_46_0/B dadda_fa_7_45_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_94_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3202 U$$3202/A U$$3224/B VGND VGND VPWR VPWR U$$3202/X sky130_fd_sc_hd__xor2_1
XU$$3213 U$$3624/A1 U$$3243/A2 _580_/Q U$$3243/B2 VGND VGND VPWR VPWR U$$3214/A sky130_fd_sc_hd__a22o_1
XFILLER_24_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3224 U$$3224/A U$$3224/B VGND VGND VPWR VPWR U$$3224/X sky130_fd_sc_hd__xor2_1
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3235 U$$632/A1 U$$3155/X U$$771/A1 U$$3156/X VGND VGND VPWR VPWR U$$3236/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$17 _441_/Q _313_/Q VGND VGND VPWR VPWR final_adder.U$$145/B1 final_adder.U$$639/A
+ sky130_fd_sc_hd__ha_1
XU$$2501 U$$2501/A U$$2533/B VGND VGND VPWR VPWR U$$2501/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$28 _452_/Q _324_/Q VGND VGND VPWR VPWR final_adder.U$$523/B1 final_adder.U$$650/A
+ sky130_fd_sc_hd__ha_1
XU$$3246 U$$3246/A U$$3270/B VGND VGND VPWR VPWR U$$3246/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2512 U$$4291/B1 U$$2534/A2 U$$4156/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2513/A
+ sky130_fd_sc_hd__a22o_1
XU$$3257 _601_/Q U$$3155/X _602_/Q U$$3156/X VGND VGND VPWR VPWR U$$3258/A sky130_fd_sc_hd__a22o_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$39 _463_/Q _335_/Q VGND VGND VPWR VPWR final_adder.U$$167/B1 final_adder.U$$661/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_104_2 dadda_fa_4_104_2/A dadda_fa_4_104_2/B dadda_fa_4_104_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/CIN dadda_fa_5_104_1/CIN sky130_fd_sc_hd__fa_2
XU$$3268 U$$3268/A U$$3270/B VGND VGND VPWR VPWR U$$3268/X sky130_fd_sc_hd__xor2_1
XU$$2523 U$$2523/A U$$2585/B VGND VGND VPWR VPWR U$$2523/X sky130_fd_sc_hd__xor2_1
XU$$3279 U$$539/A1 U$$3155/X _613_/Q U$$3156/X VGND VGND VPWR VPWR U$$3280/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2534 U$$68/A1 U$$2534/A2 U$$68/B1 U$$2534/B2 VGND VGND VPWR VPWR U$$2535/A sky130_fd_sc_hd__a22o_1
XU$$2545 U$$2545/A U$$2585/B VGND VGND VPWR VPWR U$$2545/X sky130_fd_sc_hd__xor2_1
XU$$1800 U$$1800/A U$$1918/A VGND VGND VPWR VPWR U$$1800/X sky130_fd_sc_hd__xor2_1
XU$$2556 _593_/Q U$$2470/X _594_/Q U$$2471/X VGND VGND VPWR VPWR U$$2557/A sky130_fd_sc_hd__a22o_1
XU$$1811 U$$28/B1 U$$1867/A2 U$$30/B1 U$$1867/B2 VGND VGND VPWR VPWR U$$1812/A sky130_fd_sc_hd__a22o_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1822 U$$1822/A U$$1872/B VGND VGND VPWR VPWR U$$1822/X sky130_fd_sc_hd__xor2_1
XU$$2567 U$$2567/A U$$2603/A VGND VGND VPWR VPWR U$$2567/X sky130_fd_sc_hd__xor2_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2578 U$$934/A1 U$$2470/X U$$936/A1 U$$2471/X VGND VGND VPWR VPWR U$$2579/A sky130_fd_sc_hd__a22o_1
XU$$1833 U$$2790/B1 U$$1897/A2 U$$876/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1834/A
+ sky130_fd_sc_hd__a22o_1
XU$$1844 U$$1844/A U$$1856/B VGND VGND VPWR VPWR U$$1844/X sky130_fd_sc_hd__xor2_1
XU$$2589 U$$2589/A _653_/Q VGND VGND VPWR VPWR U$$2589/X sky130_fd_sc_hd__xor2_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1855 U$$74/A1 U$$1903/A2 U$$2953/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1856/A sky130_fd_sc_hd__a22o_1
XFILLER_159_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$1866 U$$1866/A U$$1918/A VGND VGND VPWR VPWR U$$1866/X sky130_fd_sc_hd__xor2_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1877 U$$96/A1 U$$1903/A2 U$$96/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1878/A sky130_fd_sc_hd__a22o_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1888 U$$1888/A _643_/Q VGND VGND VPWR VPWR U$$1888/X sky130_fd_sc_hd__xor2_1
XU$$1899 U$$940/A1 U$$1785/X U$$942/A1 U$$1786/X VGND VGND VPWR VPWR U$$1900/A sky130_fd_sc_hd__a22o_1
XFILLER_175_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_118_0 dadda_fa_7_118_0/A dadda_fa_7_118_0/B dadda_fa_7_118_0/CIN VGND
+ VGND VPWR VPWR _543_/D _414_/D sky130_fd_sc_hd__fa_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_70_1 dadda_fa_2_70_1/A dadda_fa_2_70_1/B dadda_fa_2_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/CIN dadda_fa_3_70_2/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_63_0 dadda_fa_2_63_0/A dadda_fa_2_63_0/B dadda_fa_2_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/B dadda_fa_3_63_2/B sky130_fd_sc_hd__fa_1
Xrepeater700 _578_/Q VGND VGND VPWR VPWR U$$4170/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$507 final_adder.U$$634/A final_adder.U$$634/B final_adder.U$$507/B1
+ VGND VGND VPWR VPWR final_adder.U$$635/B sky130_fd_sc_hd__a21o_1
Xrepeater711 U$$52/A1 VGND VGND VPWR VPWR U$$50/B1 sky130_fd_sc_hd__buf_12
XFILLER_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater722 U$$3876/B1 VGND VGND VPWR VPWR U$$4289/A1 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$529 final_adder.U$$656/A final_adder.U$$656/B final_adder.U$$529/B1
+ VGND VGND VPWR VPWR final_adder.U$$657/B sky130_fd_sc_hd__a21o_1
Xrepeater733 _564_/Q VGND VGND VPWR VPWR U$$30/B1 sky130_fd_sc_hd__buf_12
Xrepeater744 _559_/Q VGND VGND VPWR VPWR U$$22/A1 sky130_fd_sc_hd__buf_12
Xrepeater755 U$$12/A1 VGND VGND VPWR VPWR U$$971/A1 sky130_fd_sc_hd__buf_12
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4470 U$$771/A1 U$$4388/X U$$771/B1 U$$4389/X VGND VGND VPWR VPWR U$$4471/A sky130_fd_sc_hd__a22o_1
XU$$4481 U$$4481/A U$$4481/B VGND VGND VPWR VPWR U$$4481/X sky130_fd_sc_hd__xor2_2
XU$$4492 U$$4492/A1 U$$4388/X U$$4494/A1 U$$4389/X VGND VGND VPWR VPWR U$$4493/A sky130_fd_sc_hd__a22o_2
XU$$3780 U$$3780/A _671_/Q VGND VGND VPWR VPWR U$$3780/X sky130_fd_sc_hd__xor2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_743__795 VGND VGND VPWR VPWR _743__795/HI U$$3011/B1 sky130_fd_sc_hd__conb_1
XFILLER_80_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3791 U$$4476/A1 U$$3795/A2 _595_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3792/A sky130_fd_sc_hd__a22o_1
XFILLER_25_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_92_2 dadda_fa_4_92_2/A dadda_fa_4_92_2/B dadda_fa_4_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/CIN dadda_fa_5_92_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_85_1 dadda_fa_4_85_1/A dadda_fa_4_85_1/B dadda_fa_4_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/B dadda_fa_5_85_1/B sky130_fd_sc_hd__fa_1
XFILLER_133_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_62_0 dadda_fa_7_62_0/A dadda_fa_7_62_0/B dadda_fa_7_62_0/CIN VGND VGND
+ VPWR VPWR _487_/D _358_/D sky130_fd_sc_hd__fa_2
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_78_0 dadda_fa_4_78_0/A dadda_fa_4_78_0/B dadda_fa_4_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/A dadda_fa_5_78_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$902 U$$902/A1 U$$928/A2 U$$902/B1 U$$928/B2 VGND VGND VPWR VPWR U$$903/A sky130_fd_sc_hd__a22o_1
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$913 U$$913/A U$$943/B VGND VGND VPWR VPWR U$$913/X sky130_fd_sc_hd__xor2_1
XU$$924 U$$924/A1 U$$928/A2 U$$926/A1 U$$928/B2 VGND VGND VPWR VPWR U$$925/A sky130_fd_sc_hd__a22o_1
XFILLER_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$935 U$$935/A U$$959/A VGND VGND VPWR VPWR U$$935/X sky130_fd_sc_hd__xor2_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$946 U$$946/A1 U$$826/X U$$948/A1 U$$827/X VGND VGND VPWR VPWR U$$947/A sky130_fd_sc_hd__a22o_1
XU$$957 U$$957/A _629_/Q VGND VGND VPWR VPWR U$$957/X sky130_fd_sc_hd__xor2_1
XU$$968 U$$968/A U$$998/B VGND VGND VPWR VPWR U$$968/X sky130_fd_sc_hd__xor2_1
XU$$1107 U$$1107/A U$$1189/B VGND VGND VPWR VPWR U$$1107/X sky130_fd_sc_hd__xor2_1
XFILLER_141_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1118 _559_/Q U$$1200/A2 U$$983/A1 U$$1200/B2 VGND VGND VPWR VPWR U$$1119/A sky130_fd_sc_hd__a22o_1
XU$$979 U$$979/A1 U$$999/A2 U$$979/B1 U$$987/B2 VGND VGND VPWR VPWR U$$980/A sky130_fd_sc_hd__a22o_1
XU$$1129 U$$1129/A U$$1189/B VGND VGND VPWR VPWR U$$1129/X sky130_fd_sc_hd__xor2_1
XFILLER_44_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_692__912 VGND VGND VPWR VPWR _692__912/HI _692__912/LO sky130_fd_sc_hd__conb_1
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_80_0 dadda_fa_3_80_0/A dadda_fa_3_80_0/B dadda_fa_3_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/B dadda_fa_4_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3010 U$$3010/A _659_/Q VGND VGND VPWR VPWR U$$3010/X sky130_fd_sc_hd__xor2_1
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_42_5 dadda_fa_2_42_5/A dadda_fa_2_42_5/B dadda_fa_2_42_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_2/A dadda_fa_4_42_0/A sky130_fd_sc_hd__fa_2
XU$$3021 U$$3021/A U$$3085/B VGND VGND VPWR VPWR U$$3021/X sky130_fd_sc_hd__xor2_1
X_727__779 VGND VGND VPWR VPWR _727__779/HI U$$2052/B1 sky130_fd_sc_hd__conb_1
XU$$3032 U$$975/B1 U$$3090/A2 U$$979/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3033/A sky130_fd_sc_hd__a22o_1
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3043 U$$3043/A U$$3129/B VGND VGND VPWR VPWR U$$3043/X sky130_fd_sc_hd__xor2_1
XU$$3054 U$$4424/A1 U$$3090/A2 U$$4289/A1 U$$3090/B2 VGND VGND VPWR VPWR U$$3055/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_35_4 U$$1939/X U$$2072/X U$$2205/X VGND VGND VPWR VPWR dadda_fa_3_36_1/CIN
+ dadda_fa_3_35_3/CIN sky130_fd_sc_hd__fa_2
XU$$2320 _612_/Q U$$2326/A2 _613_/Q U$$2326/B2 VGND VGND VPWR VPWR U$$2321/A sky130_fd_sc_hd__a22o_1
XFILLER_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$3065 U$$3065/A U$$3129/B VGND VGND VPWR VPWR U$$3065/X sky130_fd_sc_hd__xor2_1
XU$$3076 U$$3624/A1 U$$3018/X _580_/Q U$$3019/X VGND VGND VPWR VPWR U$$3077/A sky130_fd_sc_hd__a22o_1
XU$$2331 U$$2464/B VGND VGND VPWR VPWR U$$2331/Y sky130_fd_sc_hd__inv_1
XU$$3087 U$$3087/A U$$3109/B VGND VGND VPWR VPWR U$$3087/X sky130_fd_sc_hd__xor2_1
XU$$2342 U$$2342/A U$$2432/B VGND VGND VPWR VPWR U$$2342/X sky130_fd_sc_hd__xor2_1
XU$$3098 _590_/Q U$$3018/X _591_/Q U$$3019/X VGND VGND VPWR VPWR U$$3099/A sky130_fd_sc_hd__a22o_1
XU$$2353 U$$4271/A1 U$$2421/A2 U$$4273/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2354/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$2364 U$$2364/A U$$2432/B VGND VGND VPWR VPWR U$$2364/X sky130_fd_sc_hd__xor2_1
XU$$2375 U$$4291/B1 U$$2421/A2 U$$48/A1 U$$2421/B2 VGND VGND VPWR VPWR U$$2376/A sky130_fd_sc_hd__a22o_1
XU$$1630 U$$1630/A _639_/Q VGND VGND VPWR VPWR U$$1630/X sky130_fd_sc_hd__xor2_1
XFILLER_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1641 U$$956/A1 U$$1641/A2 U$$1641/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1642/A
+ sky130_fd_sc_hd__a22o_1
XU$$2386 U$$2386/A U$$2436/B VGND VGND VPWR VPWR U$$2386/X sky130_fd_sc_hd__xor2_1
XU$$2397 _582_/Q U$$2333/X U$$70/A1 U$$2334/X VGND VGND VPWR VPWR U$$2398/A sky130_fd_sc_hd__a22o_1
XU$$1652 U$$8/A1 U$$1734/A2 U$$8/B1 U$$1734/B2 VGND VGND VPWR VPWR U$$1653/A sky130_fd_sc_hd__a22o_1
XU$$1663 U$$1663/A U$$1781/A VGND VGND VPWR VPWR U$$1663/X sky130_fd_sc_hd__xor2_1
XU$$1674 U$$30/A1 U$$1726/A2 U$$30/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1675/A sky130_fd_sc_hd__a22o_1
XU$$1685 U$$1685/A U$$1727/B VGND VGND VPWR VPWR U$$1685/X sky130_fd_sc_hd__xor2_1
XU$$1696 U$$50/B1 U$$1726/A2 U$$876/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1697/A sky130_fd_sc_hd__a22o_1
XFILLER_175_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_95_0 dadda_fa_5_95_0/A dadda_fa_5_95_0/B dadda_fa_5_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/A dadda_fa_6_95_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$304 final_adder.U$$304/A final_adder.U$$304/B VGND VGND VPWR VPWR
+ final_adder.U$$344/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$315 final_adder.U$$314/A final_adder.U$$245/X final_adder.U$$247/X
+ VGND VGND VPWR VPWR final_adder.U$$315/X sky130_fd_sc_hd__a21o_1
XFILLER_97_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfinal_adder.U$$326 final_adder.U$$326/A final_adder.U$$326/B VGND VGND VPWR VPWR
+ final_adder.U$$354/A sky130_fd_sc_hd__and2_1
Xrepeater530 _669_/Q VGND VGND VPWR VPWR U$$3698/A sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$337 final_adder.U$$336/A final_adder.U$$289/X final_adder.U$$291/X
+ VGND VGND VPWR VPWR final_adder.U$$337/X sky130_fd_sc_hd__a21o_1
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater541 _663_/Q VGND VGND VPWR VPWR U$$3270/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$348 final_adder.U$$348/A final_adder.U$$348/B VGND VGND VPWR VPWR
+ final_adder.U$$348/X sky130_fd_sc_hd__and2_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater552 U$$2698/B VGND VGND VPWR VPWR U$$2694/B sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$359 final_adder.U$$358/A final_adder.U$$333/X final_adder.U$$335/X
+ VGND VGND VPWR VPWR final_adder.U$$359/X sky130_fd_sc_hd__a21o_2
Xrepeater563 _649_/Q VGND VGND VPWR VPWR U$$2327/B sky130_fd_sc_hd__buf_12
Xrepeater574 _643_/Q VGND VGND VPWR VPWR U$$1904/B sky130_fd_sc_hd__buf_12
XU$$209 U$$72/A1 U$$141/X U$$74/A1 U$$142/X VGND VGND VPWR VPWR U$$210/A sky130_fd_sc_hd__a22o_1
XFILLER_38_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater585 _635_/Q VGND VGND VPWR VPWR U$$1342/B sky130_fd_sc_hd__buf_12
Xrepeater596 _629_/Q VGND VGND VPWR VPWR U$$959/A sky130_fd_sc_hd__buf_12
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_3_111_2 U$$4086/X U$$4219/X U$$4352/X VGND VGND VPWR VPWR dadda_fa_4_112_1/CIN
+ dadda_fa_4_111_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_104_1 U$$4205/X U$$4338/X U$$4471/X VGND VGND VPWR VPWR dadda_fa_4_105_0/CIN
+ dadda_fa_4_104_2/A sky130_fd_sc_hd__fa_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_6_125_0 input157/X dadda_fa_6_125_0/B dadda_fa_6_125_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_126_0/B dadda_fa_7_125_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_0_68_4 U$$1872/X U$$2005/X U$$2138/X VGND VGND VPWR VPWR dadda_fa_1_69_7/A
+ dadda_fa_1_68_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_45_3 dadda_fa_3_45_3/A dadda_fa_3_45_3/B dadda_fa_3_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/B dadda_fa_4_45_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$710 U$$710/A U$$784/B VGND VGND VPWR VPWR U$$710/X sky130_fd_sc_hd__xor2_1
X_664_ _667_/CLK _664_/D VGND VGND VPWR VPWR _664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_38_2 dadda_fa_3_38_2/A dadda_fa_3_38_2/B dadda_fa_3_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/A dadda_fa_4_38_2/B sky130_fd_sc_hd__fa_1
XFILLER_17_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$721 U$$36/A1 U$$785/A2 U$$38/A1 U$$785/B2 VGND VGND VPWR VPWR U$$722/A sky130_fd_sc_hd__a22o_1
XU$$732 U$$732/A U$$784/B VGND VGND VPWR VPWR U$$732/X sky130_fd_sc_hd__xor2_1
XU$$743 U$$880/A1 U$$785/A2 U$$60/A1 U$$785/B2 VGND VGND VPWR VPWR U$$744/A sky130_fd_sc_hd__a22o_1
XU$$754 U$$754/A U$$784/B VGND VGND VPWR VPWR U$$754/X sky130_fd_sc_hd__xor2_1
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XU$$765 U$$765/A1 U$$689/X U$$82/A1 U$$690/X VGND VGND VPWR VPWR U$$766/A sky130_fd_sc_hd__a22o_1
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_595_ _595_/CLK _595_/D VGND VGND VPWR VPWR _595_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$776 U$$776/A _627_/Q VGND VGND VPWR VPWR U$$776/X sky130_fd_sc_hd__xor2_1
XU$$787 U$$924/A1 U$$817/A2 U$$787/B1 U$$817/B2 VGND VGND VPWR VPWR U$$788/A sky130_fd_sc_hd__a22o_1
XU$$798 U$$798/A U$$822/A VGND VGND VPWR VPWR U$$798/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_2_27_2 U$$859/X U$$992/X VGND VGND VPWR VPWR dadda_fa_3_28_2/CIN dadda_fa_4_27_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_2_40_2 U$$2348/X U$$2481/X U$$2614/X VGND VGND VPWR VPWR dadda_fa_3_41_1/A
+ dadda_fa_3_40_3/A sky130_fd_sc_hd__fa_1
XFILLER_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_33_1 U$$472/X U$$605/X U$$738/X VGND VGND VPWR VPWR dadda_fa_3_34_0/CIN
+ dadda_fa_3_33_2/CIN sky130_fd_sc_hd__fa_2
XU$$2150 U$$2150/A _647_/Q VGND VGND VPWR VPWR U$$2150/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_10_0 U$$692/X U$$784/B input140/X VGND VGND VPWR VPWR dadda_fa_6_11_0/A
+ dadda_fa_6_10_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_26_0 U$$59/X U$$192/X U$$325/X VGND VGND VPWR VPWR dadda_fa_3_27_2/B dadda_fa_3_26_3/B
+ sky130_fd_sc_hd__fa_2
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2161 U$$654/A1 U$$2161/A2 U$$930/A1 U$$2161/B2 VGND VGND VPWR VPWR U$$2162/A sky130_fd_sc_hd__a22o_1
XU$$2172 U$$2172/A U$$2186/B VGND VGND VPWR VPWR U$$2172/X sky130_fd_sc_hd__xor2_1
XU$$2183 U$$950/A1 U$$2189/A2 U$$952/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2184/A sky130_fd_sc_hd__a22o_1
XFILLER_179_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2194 _649_/Q VGND VGND VPWR VPWR U$$2194/Y sky130_fd_sc_hd__inv_1
XU$$1460 U$$912/A1 U$$1472/A2 U$$92/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1461/A sky130_fd_sc_hd__a22o_1
XU$$1471 U$$1471/A U$$1505/B VGND VGND VPWR VPWR U$$1471/X sky130_fd_sc_hd__xor2_1
XU$$1482 _604_/Q U$$1374/X U$$799/A1 U$$1375/X VGND VGND VPWR VPWR U$$1483/A sky130_fd_sc_hd__a22o_1
XU$$1493 U$$1493/A U$$1505/B VGND VGND VPWR VPWR U$$1493/X sky130_fd_sc_hd__xor2_1
XFILLER_176_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_85_4 U$$3103/X U$$3236/X U$$3369/X VGND VGND VPWR VPWR dadda_fa_2_86_3/CIN
+ dadda_fa_2_85_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_1_78_3 U$$2424/X U$$2557/X U$$2690/X VGND VGND VPWR VPWR dadda_fa_2_79_1/B
+ dadda_fa_2_78_4/B sky130_fd_sc_hd__fa_1
XFILLER_44_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_55_2 dadda_fa_4_55_2/A dadda_fa_4_55_2/B dadda_fa_4_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/CIN dadda_fa_5_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$101 _525_/Q _397_/Q VGND VGND VPWR VPWR final_adder.U$$229/B1 final_adder.U$$723/A
+ sky130_fd_sc_hd__ha_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$112 _536_/Q _408_/Q VGND VGND VPWR VPWR final_adder.U$$607/B1 final_adder.U$$734/A
+ sky130_fd_sc_hd__ha_1
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$123 _547_/Q _419_/Q VGND VGND VPWR VPWR final_adder.U$$251/B1 final_adder.U$$745/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_4_48_1 dadda_fa_4_48_1/A dadda_fa_4_48_1/B dadda_fa_4_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/B dadda_fa_5_48_1/B sky130_fd_sc_hd__fa_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$134 final_adder.U$$7/SUM final_adder.U$$628/A VGND VGND VPWR VPWR
+ final_adder.U$$258/A sky130_fd_sc_hd__and2_1
XFILLER_181_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$145 final_adder.U$$639/A final_adder.U$$511/B1 final_adder.U$$145/B1
+ VGND VGND VPWR VPWR final_adder.U$$145/X sky130_fd_sc_hd__a21o_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_25_0 dadda_fa_7_25_0/A dadda_fa_7_25_0/B dadda_fa_7_25_0/CIN VGND VGND
+ VPWR VPWR _450_/D _321_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$156 final_adder.U$$651/A final_adder.U$$650/A VGND VGND VPWR VPWR
+ final_adder.U$$270/B sky130_fd_sc_hd__and2_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$167 final_adder.U$$661/A final_adder.U$$533/B1 final_adder.U$$167/B1
+ VGND VGND VPWR VPWR final_adder.U$$167/X sky130_fd_sc_hd__a21o_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$178 final_adder.U$$673/A final_adder.U$$672/A VGND VGND VPWR VPWR
+ final_adder.U$$280/A sky130_fd_sc_hd__and2_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$189 final_adder.U$$683/A final_adder.U$$555/B1 final_adder.U$$189/B1
+ VGND VGND VPWR VPWR final_adder.U$$189/X sky130_fd_sc_hd__a21o_1
Xrepeater393 U$$4381/A2 VGND VGND VPWR VPWR U$$4377/A2 sky130_fd_sc_hd__buf_12
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_380_ _510_/CLK _380_/D VGND VGND VPWR VPWR _380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_73_2 U$$1483/X U$$1616/X U$$1749/X VGND VGND VPWR VPWR dadda_fa_1_74_8/A
+ dadda_fa_2_73_0/A sky130_fd_sc_hd__fa_2
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput130 c[100] VGND VGND VPWR VPWR input130/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput141 c[110] VGND VGND VPWR VPWR input141/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_50_1 dadda_fa_3_50_1/A dadda_fa_3_50_1/B dadda_fa_3_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/CIN dadda_fa_4_50_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_0_66_1 U$$538/X U$$671/X U$$804/X VGND VGND VPWR VPWR dadda_fa_1_67_5/CIN
+ dadda_fa_1_66_7/CIN sky130_fd_sc_hd__fa_1
Xinput152 c[120] VGND VGND VPWR VPWR input152/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 c[15] VGND VGND VPWR VPWR input163/X sky130_fd_sc_hd__clkbuf_2
Xinput174 c[25] VGND VGND VPWR VPWR input174/X sky130_fd_sc_hd__buf_2
XFILLER_110_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_43_0 dadda_fa_3_43_0/A dadda_fa_3_43_0/B dadda_fa_3_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/B dadda_fa_4_43_1/CIN sky130_fd_sc_hd__fa_1
Xinput185 c[35] VGND VGND VPWR VPWR input185/X sky130_fd_sc_hd__buf_4
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput196 c[45] VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_59_0 U$$125/X U$$258/X U$$391/X VGND VGND VPWR VPWR dadda_fa_1_60_6/B
+ dadda_fa_1_59_8/A sky130_fd_sc_hd__fa_1
XFILLER_91_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$690 final_adder.U$$690/A final_adder.U$$690/B VGND VGND VPWR VPWR
+ _236_/D sky130_fd_sc_hd__xor2_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$540 U$$540/A _623_/Q VGND VGND VPWR VPWR U$$540/X sky130_fd_sc_hd__xor2_1
X_647_ _647_/CLK _647_/D VGND VGND VPWR VPWR _647_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$551 _625_/Q U$$551/B VGND VGND VPWR VPWR U$$551/X sky130_fd_sc_hd__and2_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$562 U$$12/B1 U$$682/A2 U$$16/A1 U$$553/X VGND VGND VPWR VPWR U$$563/A sky130_fd_sc_hd__a22o_1
XU$$573 U$$573/A U$$623/B VGND VGND VPWR VPWR U$$573/X sky130_fd_sc_hd__xor2_1
XFILLER_189_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$584 U$$36/A1 U$$626/A2 U$$38/A1 U$$553/X VGND VGND VPWR VPWR U$$585/A sky130_fd_sc_hd__a22o_1
XFILLER_189_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$595 U$$595/A U$$623/B VGND VGND VPWR VPWR U$$595/X sky130_fd_sc_hd__xor2_1
X_578_ _578_/CLK _578_/D VGND VGND VPWR VPWR _578_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_100_0 dadda_fa_7_100_0/A dadda_fa_7_100_0/B dadda_fa_7_100_0/CIN VGND
+ VGND VPWR VPWR _525_/D _396_/D sky130_fd_sc_hd__fa_2
XFILLER_173_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_95_3 U$$3788/X U$$3921/X U$$4054/X VGND VGND VPWR VPWR dadda_fa_3_96_1/B
+ dadda_fa_3_95_3/B sky130_fd_sc_hd__fa_1
XFILLER_160_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_88_2 U$$4306/X U$$4439/X input243/X VGND VGND VPWR VPWR dadda_fa_3_89_1/A
+ dadda_fa_3_88_3/A sky130_fd_sc_hd__fa_2
XFILLER_113_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xdadda_fa_5_65_1 dadda_fa_5_65_1/A dadda_fa_5_65_1/B dadda_fa_5_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/B dadda_fa_7_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_58_0 dadda_fa_5_58_0/A dadda_fa_5_58_0/B dadda_fa_5_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/A dadda_fa_6_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

