VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM32_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 1123.780 BY 185.440 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 125.160 1123.780 125.760 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 138.760 1123.780 139.360 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 151.680 1123.780 152.280 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 165.280 1123.780 165.880 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 178.200 1123.780 178.800 ;
    END
  END A0[4]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.000 40.080 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.000 66.600 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.000 93.120 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 2.000 119.640 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 2.000 146.160 ;
    END
  END A1[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.000 13.560 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 0.000 904.270 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 0.000 974.650 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 0.000 1062.510 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 0.000 1114.950 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 183.440 4.510 185.440 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 183.440 91.910 185.440 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 183.440 109.850 185.440 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 183.440 127.330 185.440 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 183.440 144.810 185.440 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 183.440 162.290 185.440 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 183.440 179.770 185.440 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 183.440 197.250 185.440 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 183.440 215.190 185.440 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 183.440 232.670 185.440 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 183.440 250.150 185.440 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 183.440 13.250 185.440 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 183.440 267.630 185.440 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 183.440 276.370 185.440 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 183.440 285.110 185.440 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 183.440 293.850 185.440 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 183.440 302.590 185.440 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 183.440 311.790 185.440 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 183.440 320.530 185.440 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 183.440 329.270 185.440 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 183.440 338.010 185.440 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 183.440 346.750 185.440 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 183.440 21.990 185.440 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 183.440 355.490 185.440 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 183.440 364.230 185.440 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 183.440 372.970 185.440 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 183.440 381.710 185.440 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 183.440 390.450 185.440 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 183.440 399.190 185.440 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 183.440 407.930 185.440 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 183.440 417.130 185.440 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 183.440 425.870 185.440 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 183.440 434.610 185.440 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 183.440 30.730 185.440 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 183.440 443.350 185.440 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 183.440 452.090 185.440 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 183.440 460.830 185.440 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 183.440 469.570 185.440 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 183.440 478.310 185.440 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 183.440 487.050 185.440 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 183.440 495.790 185.440 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 183.440 504.530 185.440 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 183.440 513.270 185.440 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 183.440 522.470 185.440 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 183.440 39.470 185.440 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 183.440 531.210 185.440 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 183.440 539.950 185.440 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 183.440 548.690 185.440 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 183.440 557.430 185.440 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 183.440 566.170 185.440 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 183.440 574.910 185.440 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 183.440 583.650 185.440 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 183.440 592.390 185.440 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 183.440 601.130 185.440 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 183.440 609.870 185.440 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 183.440 48.210 185.440 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 183.440 619.070 185.440 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 183.440 627.810 185.440 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 183.440 636.550 185.440 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 183.440 645.290 185.440 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 183.440 56.950 185.440 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 183.440 65.690 185.440 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 183.440 74.430 185.440 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 183.440 83.170 185.440 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 183.440 100.650 185.440 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 183.440 654.030 185.440 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 183.440 662.770 185.440 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 183.440 671.510 185.440 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 183.440 680.250 185.440 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 183.440 688.990 185.440 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 183.440 697.730 185.440 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 183.440 706.470 185.440 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 183.440 715.210 185.440 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 183.440 724.410 185.440 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 183.440 733.150 185.440 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 183.440 118.590 185.440 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 183.440 741.890 185.440 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 183.440 750.630 185.440 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 183.440 759.370 185.440 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 183.440 768.110 185.440 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 183.440 776.850 185.440 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 183.440 785.590 185.440 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 183.440 794.330 185.440 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 183.440 803.070 185.440 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 183.440 811.810 185.440 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 183.440 820.550 185.440 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 183.440 136.070 185.440 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 183.440 829.750 185.440 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 183.440 838.490 185.440 ;
    END
  END Do1[31]
  PIN Do1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 183.440 847.230 185.440 ;
    END
  END Do1[32]
  PIN Do1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 183.440 855.970 185.440 ;
    END
  END Do1[33]
  PIN Do1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 183.440 864.710 185.440 ;
    END
  END Do1[34]
  PIN Do1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 183.440 873.450 185.440 ;
    END
  END Do1[35]
  PIN Do1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 183.440 882.190 185.440 ;
    END
  END Do1[36]
  PIN Do1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 183.440 890.930 185.440 ;
    END
  END Do1[37]
  PIN Do1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 183.440 899.670 185.440 ;
    END
  END Do1[38]
  PIN Do1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 183.440 908.410 185.440 ;
    END
  END Do1[39]
  PIN Do1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 183.440 153.550 185.440 ;
    END
  END Do1[3]
  PIN Do1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 183.440 917.150 185.440 ;
    END
  END Do1[40]
  PIN Do1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 183.440 926.350 185.440 ;
    END
  END Do1[41]
  PIN Do1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 183.440 935.090 185.440 ;
    END
  END Do1[42]
  PIN Do1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 183.440 943.830 185.440 ;
    END
  END Do1[43]
  PIN Do1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 183.440 952.570 185.440 ;
    END
  END Do1[44]
  PIN Do1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 183.440 961.310 185.440 ;
    END
  END Do1[45]
  PIN Do1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 183.440 970.050 185.440 ;
    END
  END Do1[46]
  PIN Do1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 183.440 978.790 185.440 ;
    END
  END Do1[47]
  PIN Do1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 183.440 987.530 185.440 ;
    END
  END Do1[48]
  PIN Do1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 183.440 996.270 185.440 ;
    END
  END Do1[49]
  PIN Do1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 183.440 171.030 185.440 ;
    END
  END Do1[4]
  PIN Do1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 183.440 1005.010 185.440 ;
    END
  END Do1[50]
  PIN Do1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.470 183.440 1013.750 185.440 ;
    END
  END Do1[51]
  PIN Do1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 183.440 1022.490 185.440 ;
    END
  END Do1[52]
  PIN Do1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 183.440 1031.690 185.440 ;
    END
  END Do1[53]
  PIN Do1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 183.440 1040.430 185.440 ;
    END
  END Do1[54]
  PIN Do1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 183.440 1049.170 185.440 ;
    END
  END Do1[55]
  PIN Do1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.630 183.440 1057.910 185.440 ;
    END
  END Do1[56]
  PIN Do1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 183.440 1066.650 185.440 ;
    END
  END Do1[57]
  PIN Do1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 183.440 1075.390 185.440 ;
    END
  END Do1[58]
  PIN Do1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 183.440 1084.130 185.440 ;
    END
  END Do1[59]
  PIN Do1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 183.440 188.510 185.440 ;
    END
  END Do1[5]
  PIN Do1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 183.440 1092.870 185.440 ;
    END
  END Do1[60]
  PIN Do1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 183.440 1101.610 185.440 ;
    END
  END Do1[61]
  PIN Do1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 183.440 1110.350 185.440 ;
    END
  END Do1[62]
  PIN Do1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 183.440 1119.090 185.440 ;
    END
  END Do1[63]
  PIN Do1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 183.440 205.990 185.440 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 183.440 223.930 185.440 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 183.440 241.410 185.440 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 183.440 258.890 185.440 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 6.160 1123.780 6.760 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 2.000 172.680 ;
    END
  END EN1
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.210 2.480 99.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.210 2.480 279.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.210 2.480 459.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.210 2.480 639.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.210 2.480 819.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.210 2.480 999.310 182.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.210 2.480 9.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.210 2.480 189.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.210 2.480 369.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.210 2.480 549.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.210 2.480 729.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.210 2.480 909.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1086.210 2.480 1089.310 182.480 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 19.080 1123.780 19.680 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 32.680 1123.780 33.280 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 45.600 1123.780 46.200 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 59.200 1123.780 59.800 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 72.120 1123.780 72.720 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 85.720 1123.780 86.320 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 98.640 1123.780 99.240 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1121.780 112.240 1123.780 112.840 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 1121.020 98.005 ;
      LAYER met1 ;
        RECT 0.990 0.380 1121.020 184.240 ;
      LAYER met2 ;
        RECT 1.020 183.160 3.950 184.270 ;
        RECT 4.790 183.160 12.690 184.270 ;
        RECT 13.530 183.160 21.430 184.270 ;
        RECT 22.270 183.160 30.170 184.270 ;
        RECT 31.010 183.160 38.910 184.270 ;
        RECT 39.750 183.160 47.650 184.270 ;
        RECT 48.490 183.160 56.390 184.270 ;
        RECT 57.230 183.160 65.130 184.270 ;
        RECT 65.970 183.160 73.870 184.270 ;
        RECT 74.710 183.160 82.610 184.270 ;
        RECT 83.450 183.160 91.350 184.270 ;
        RECT 92.190 183.160 100.090 184.270 ;
        RECT 100.930 183.160 109.290 184.270 ;
        RECT 110.130 183.160 118.030 184.270 ;
        RECT 118.870 183.160 126.770 184.270 ;
        RECT 127.610 183.160 135.510 184.270 ;
        RECT 136.350 183.160 144.250 184.270 ;
        RECT 145.090 183.160 152.990 184.270 ;
        RECT 153.830 183.160 161.730 184.270 ;
        RECT 162.570 183.160 170.470 184.270 ;
        RECT 171.310 183.160 179.210 184.270 ;
        RECT 180.050 183.160 187.950 184.270 ;
        RECT 188.790 183.160 196.690 184.270 ;
        RECT 197.530 183.160 205.430 184.270 ;
        RECT 206.270 183.160 214.630 184.270 ;
        RECT 215.470 183.160 223.370 184.270 ;
        RECT 224.210 183.160 232.110 184.270 ;
        RECT 232.950 183.160 240.850 184.270 ;
        RECT 241.690 183.160 249.590 184.270 ;
        RECT 250.430 183.160 258.330 184.270 ;
        RECT 259.170 183.160 267.070 184.270 ;
        RECT 267.910 183.160 275.810 184.270 ;
        RECT 276.650 183.160 284.550 184.270 ;
        RECT 285.390 183.160 293.290 184.270 ;
        RECT 294.130 183.160 302.030 184.270 ;
        RECT 302.870 183.160 311.230 184.270 ;
        RECT 312.070 183.160 319.970 184.270 ;
        RECT 320.810 183.160 328.710 184.270 ;
        RECT 329.550 183.160 337.450 184.270 ;
        RECT 338.290 183.160 346.190 184.270 ;
        RECT 347.030 183.160 354.930 184.270 ;
        RECT 355.770 183.160 363.670 184.270 ;
        RECT 364.510 183.160 372.410 184.270 ;
        RECT 373.250 183.160 381.150 184.270 ;
        RECT 381.990 183.160 389.890 184.270 ;
        RECT 390.730 183.160 398.630 184.270 ;
        RECT 399.470 183.160 407.370 184.270 ;
        RECT 408.210 183.160 416.570 184.270 ;
        RECT 417.410 183.160 425.310 184.270 ;
        RECT 426.150 183.160 434.050 184.270 ;
        RECT 434.890 183.160 442.790 184.270 ;
        RECT 443.630 183.160 451.530 184.270 ;
        RECT 452.370 183.160 460.270 184.270 ;
        RECT 461.110 183.160 469.010 184.270 ;
        RECT 469.850 183.160 477.750 184.270 ;
        RECT 478.590 183.160 486.490 184.270 ;
        RECT 487.330 183.160 495.230 184.270 ;
        RECT 496.070 183.160 503.970 184.270 ;
        RECT 504.810 183.160 512.710 184.270 ;
        RECT 513.550 183.160 521.910 184.270 ;
        RECT 522.750 183.160 530.650 184.270 ;
        RECT 531.490 183.160 539.390 184.270 ;
        RECT 540.230 183.160 548.130 184.270 ;
        RECT 548.970 183.160 556.870 184.270 ;
        RECT 557.710 183.160 565.610 184.270 ;
        RECT 566.450 183.160 574.350 184.270 ;
        RECT 575.190 183.160 583.090 184.270 ;
        RECT 583.930 183.160 591.830 184.270 ;
        RECT 592.670 183.160 600.570 184.270 ;
        RECT 601.410 183.160 609.310 184.270 ;
        RECT 610.150 183.160 618.510 184.270 ;
        RECT 619.350 183.160 627.250 184.270 ;
        RECT 628.090 183.160 635.990 184.270 ;
        RECT 636.830 183.160 644.730 184.270 ;
        RECT 645.570 183.160 653.470 184.270 ;
        RECT 654.310 183.160 662.210 184.270 ;
        RECT 663.050 183.160 670.950 184.270 ;
        RECT 671.790 183.160 679.690 184.270 ;
        RECT 680.530 183.160 688.430 184.270 ;
        RECT 689.270 183.160 697.170 184.270 ;
        RECT 698.010 183.160 705.910 184.270 ;
        RECT 706.750 183.160 714.650 184.270 ;
        RECT 715.490 183.160 723.850 184.270 ;
        RECT 724.690 183.160 732.590 184.270 ;
        RECT 733.430 183.160 741.330 184.270 ;
        RECT 742.170 183.160 750.070 184.270 ;
        RECT 750.910 183.160 758.810 184.270 ;
        RECT 759.650 183.160 767.550 184.270 ;
        RECT 768.390 183.160 776.290 184.270 ;
        RECT 777.130 183.160 785.030 184.270 ;
        RECT 785.870 183.160 793.770 184.270 ;
        RECT 794.610 183.160 802.510 184.270 ;
        RECT 803.350 183.160 811.250 184.270 ;
        RECT 812.090 183.160 819.990 184.270 ;
        RECT 820.830 183.160 829.190 184.270 ;
        RECT 830.030 183.160 837.930 184.270 ;
        RECT 838.770 183.160 846.670 184.270 ;
        RECT 847.510 183.160 855.410 184.270 ;
        RECT 856.250 183.160 864.150 184.270 ;
        RECT 864.990 183.160 872.890 184.270 ;
        RECT 873.730 183.160 881.630 184.270 ;
        RECT 882.470 183.160 890.370 184.270 ;
        RECT 891.210 183.160 899.110 184.270 ;
        RECT 899.950 183.160 907.850 184.270 ;
        RECT 908.690 183.160 916.590 184.270 ;
        RECT 917.430 183.160 925.790 184.270 ;
        RECT 926.630 183.160 934.530 184.270 ;
        RECT 935.370 183.160 943.270 184.270 ;
        RECT 944.110 183.160 952.010 184.270 ;
        RECT 952.850 183.160 960.750 184.270 ;
        RECT 961.590 183.160 969.490 184.270 ;
        RECT 970.330 183.160 978.230 184.270 ;
        RECT 979.070 183.160 986.970 184.270 ;
        RECT 987.810 183.160 995.710 184.270 ;
        RECT 996.550 183.160 1004.450 184.270 ;
        RECT 1005.290 183.160 1013.190 184.270 ;
        RECT 1014.030 183.160 1021.930 184.270 ;
        RECT 1022.770 183.160 1031.130 184.270 ;
        RECT 1031.970 183.160 1039.870 184.270 ;
        RECT 1040.710 183.160 1048.610 184.270 ;
        RECT 1049.450 183.160 1057.350 184.270 ;
        RECT 1058.190 183.160 1066.090 184.270 ;
        RECT 1066.930 183.160 1074.830 184.270 ;
        RECT 1075.670 183.160 1083.570 184.270 ;
        RECT 1084.410 183.160 1092.310 184.270 ;
        RECT 1093.150 183.160 1101.050 184.270 ;
        RECT 1101.890 183.160 1109.790 184.270 ;
        RECT 1110.630 183.160 1118.530 184.270 ;
        RECT 1119.370 183.160 1120.000 184.270 ;
        RECT 1.020 2.280 1120.000 183.160 ;
        RECT 1.020 0.155 8.550 2.280 ;
        RECT 9.390 0.155 26.030 2.280 ;
        RECT 26.870 0.155 43.510 2.280 ;
        RECT 44.350 0.155 60.990 2.280 ;
        RECT 61.830 0.155 78.470 2.280 ;
        RECT 79.310 0.155 95.950 2.280 ;
        RECT 96.790 0.155 113.890 2.280 ;
        RECT 114.730 0.155 131.370 2.280 ;
        RECT 132.210 0.155 148.850 2.280 ;
        RECT 149.690 0.155 166.330 2.280 ;
        RECT 167.170 0.155 183.810 2.280 ;
        RECT 184.650 0.155 201.290 2.280 ;
        RECT 202.130 0.155 219.230 2.280 ;
        RECT 220.070 0.155 236.710 2.280 ;
        RECT 237.550 0.155 254.190 2.280 ;
        RECT 255.030 0.155 271.670 2.280 ;
        RECT 272.510 0.155 289.150 2.280 ;
        RECT 289.990 0.155 306.630 2.280 ;
        RECT 307.470 0.155 324.570 2.280 ;
        RECT 325.410 0.155 342.050 2.280 ;
        RECT 342.890 0.155 359.530 2.280 ;
        RECT 360.370 0.155 377.010 2.280 ;
        RECT 377.850 0.155 394.490 2.280 ;
        RECT 395.330 0.155 411.970 2.280 ;
        RECT 412.810 0.155 429.910 2.280 ;
        RECT 430.750 0.155 447.390 2.280 ;
        RECT 448.230 0.155 464.870 2.280 ;
        RECT 465.710 0.155 482.350 2.280 ;
        RECT 483.190 0.155 499.830 2.280 ;
        RECT 500.670 0.155 517.310 2.280 ;
        RECT 518.150 0.155 535.250 2.280 ;
        RECT 536.090 0.155 552.730 2.280 ;
        RECT 553.570 0.155 570.210 2.280 ;
        RECT 571.050 0.155 587.690 2.280 ;
        RECT 588.530 0.155 605.170 2.280 ;
        RECT 606.010 0.155 623.110 2.280 ;
        RECT 623.950 0.155 640.590 2.280 ;
        RECT 641.430 0.155 658.070 2.280 ;
        RECT 658.910 0.155 675.550 2.280 ;
        RECT 676.390 0.155 693.030 2.280 ;
        RECT 693.870 0.155 710.510 2.280 ;
        RECT 711.350 0.155 728.450 2.280 ;
        RECT 729.290 0.155 745.930 2.280 ;
        RECT 746.770 0.155 763.410 2.280 ;
        RECT 764.250 0.155 780.890 2.280 ;
        RECT 781.730 0.155 798.370 2.280 ;
        RECT 799.210 0.155 815.850 2.280 ;
        RECT 816.690 0.155 833.790 2.280 ;
        RECT 834.630 0.155 851.270 2.280 ;
        RECT 852.110 0.155 868.750 2.280 ;
        RECT 869.590 0.155 886.230 2.280 ;
        RECT 887.070 0.155 903.710 2.280 ;
        RECT 904.550 0.155 921.190 2.280 ;
        RECT 922.030 0.155 939.130 2.280 ;
        RECT 939.970 0.155 956.610 2.280 ;
        RECT 957.450 0.155 974.090 2.280 ;
        RECT 974.930 0.155 991.570 2.280 ;
        RECT 992.410 0.155 1009.050 2.280 ;
        RECT 1009.890 0.155 1026.530 2.280 ;
        RECT 1027.370 0.155 1044.470 2.280 ;
        RECT 1045.310 0.155 1061.950 2.280 ;
        RECT 1062.790 0.155 1079.430 2.280 ;
        RECT 1080.270 0.155 1096.910 2.280 ;
        RECT 1097.750 0.155 1114.390 2.280 ;
        RECT 1115.230 0.155 1120.000 2.280 ;
      LAYER met3 ;
        RECT 2.000 179.200 1121.780 182.405 ;
        RECT 2.000 177.800 1121.380 179.200 ;
        RECT 2.000 173.080 1121.780 177.800 ;
        RECT 2.400 171.680 1121.780 173.080 ;
        RECT 2.000 166.280 1121.780 171.680 ;
        RECT 2.000 164.880 1121.380 166.280 ;
        RECT 2.000 152.680 1121.780 164.880 ;
        RECT 2.000 151.280 1121.380 152.680 ;
        RECT 2.000 146.560 1121.780 151.280 ;
        RECT 2.400 145.160 1121.780 146.560 ;
        RECT 2.000 139.760 1121.780 145.160 ;
        RECT 2.000 138.360 1121.380 139.760 ;
        RECT 2.000 126.160 1121.780 138.360 ;
        RECT 2.000 124.760 1121.380 126.160 ;
        RECT 2.000 120.040 1121.780 124.760 ;
        RECT 2.400 118.640 1121.780 120.040 ;
        RECT 2.000 113.240 1121.780 118.640 ;
        RECT 2.000 111.840 1121.380 113.240 ;
        RECT 2.000 99.640 1121.780 111.840 ;
        RECT 2.000 98.240 1121.380 99.640 ;
        RECT 2.000 93.520 1121.780 98.240 ;
        RECT 2.400 92.120 1121.780 93.520 ;
        RECT 2.000 86.720 1121.780 92.120 ;
        RECT 2.000 85.320 1121.380 86.720 ;
        RECT 2.000 73.120 1121.780 85.320 ;
        RECT 2.000 71.720 1121.380 73.120 ;
        RECT 2.000 67.000 1121.780 71.720 ;
        RECT 2.400 65.600 1121.780 67.000 ;
        RECT 2.000 60.200 1121.780 65.600 ;
        RECT 2.000 58.800 1121.380 60.200 ;
        RECT 2.000 46.600 1121.780 58.800 ;
        RECT 2.000 45.200 1121.380 46.600 ;
        RECT 2.000 40.480 1121.780 45.200 ;
        RECT 2.400 39.080 1121.780 40.480 ;
        RECT 2.000 33.680 1121.780 39.080 ;
        RECT 2.000 32.280 1121.380 33.680 ;
        RECT 2.000 20.080 1121.780 32.280 ;
        RECT 2.000 18.680 1121.380 20.080 ;
        RECT 2.000 13.960 1121.780 18.680 ;
        RECT 2.400 12.560 1121.780 13.960 ;
        RECT 2.000 7.160 1121.780 12.560 ;
        RECT 2.000 5.760 1121.380 7.160 ;
        RECT 2.000 0.175 1121.780 5.760 ;
      LAYER met4 ;
        RECT 16.855 2.215 95.810 175.265 ;
        RECT 99.710 2.215 185.810 175.265 ;
        RECT 189.710 2.215 275.810 175.265 ;
        RECT 279.710 2.215 365.810 175.265 ;
        RECT 369.710 2.215 455.810 175.265 ;
        RECT 459.710 2.215 545.810 175.265 ;
        RECT 549.710 2.215 635.810 175.265 ;
        RECT 639.710 2.215 725.810 175.265 ;
        RECT 729.710 2.215 815.810 175.265 ;
        RECT 819.710 2.215 905.810 175.265 ;
        RECT 909.710 2.215 995.810 175.265 ;
        RECT 999.710 2.215 1077.025 175.265 ;
  END
END RAM32_1RW1R
END LIBRARY

