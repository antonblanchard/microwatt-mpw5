magic
tech sky130A
magscale 1 2
timestamp 1645351752
<< obsli1 >>
rect 4048 20111 314916 177361
<< obsm1 >>
rect 290 8 318674 197464
<< metal2 >>
rect 2502 197072 2558 197472
rect 7470 197072 7526 197472
rect 12438 197072 12494 197472
rect 17406 197072 17462 197472
rect 22374 197072 22430 197472
rect 27342 197072 27398 197472
rect 32402 197072 32458 197472
rect 37370 197072 37426 197472
rect 42338 197072 42394 197472
rect 47306 197072 47362 197472
rect 52274 197072 52330 197472
rect 57242 197072 57298 197472
rect 62302 197072 62358 197472
rect 67270 197072 67326 197472
rect 72238 197072 72294 197472
rect 77206 197072 77262 197472
rect 82174 197072 82230 197472
rect 87142 197072 87198 197472
rect 92202 197072 92258 197472
rect 97170 197072 97226 197472
rect 102138 197072 102194 197472
rect 107106 197072 107162 197472
rect 112074 197072 112130 197472
rect 117042 197072 117098 197472
rect 122102 197072 122158 197472
rect 127070 197072 127126 197472
rect 132038 197072 132094 197472
rect 137006 197072 137062 197472
rect 141974 197072 142030 197472
rect 146942 197072 146998 197472
rect 152002 197072 152058 197472
rect 156970 197072 157026 197472
rect 161938 197072 161994 197472
rect 166906 197072 166962 197472
rect 171874 197072 171930 197472
rect 176934 197072 176990 197472
rect 181902 197072 181958 197472
rect 186870 197072 186926 197472
rect 191838 197072 191894 197472
rect 196806 197072 196862 197472
rect 201774 197072 201830 197472
rect 206834 197072 206890 197472
rect 211802 197072 211858 197472
rect 216770 197072 216826 197472
rect 221738 197072 221794 197472
rect 226706 197072 226762 197472
rect 231674 197072 231730 197472
rect 236734 197072 236790 197472
rect 241702 197072 241758 197472
rect 246670 197072 246726 197472
rect 251638 197072 251694 197472
rect 256606 197072 256662 197472
rect 261574 197072 261630 197472
rect 266634 197072 266690 197472
rect 271602 197072 271658 197472
rect 276570 197072 276626 197472
rect 281538 197072 281594 197472
rect 286506 197072 286562 197472
rect 291474 197072 291530 197472
rect 296534 197072 296590 197472
rect 301502 197072 301558 197472
rect 306470 197072 306526 197472
rect 311438 197072 311494 197472
rect 316406 197072 316462 197472
rect 2502 0 2558 400
rect 7470 0 7526 400
rect 12438 0 12494 400
rect 17406 0 17462 400
rect 22374 0 22430 400
rect 27342 0 27398 400
rect 32402 0 32458 400
rect 37370 0 37426 400
rect 42338 0 42394 400
rect 47306 0 47362 400
rect 52274 0 52330 400
rect 57242 0 57298 400
rect 62302 0 62358 400
rect 67270 0 67326 400
rect 72238 0 72294 400
rect 77206 0 77262 400
rect 82174 0 82230 400
rect 87142 0 87198 400
rect 92202 0 92258 400
rect 97170 0 97226 400
rect 102138 0 102194 400
rect 107106 0 107162 400
rect 112074 0 112130 400
rect 117042 0 117098 400
rect 122102 0 122158 400
rect 127070 0 127126 400
rect 132038 0 132094 400
rect 137006 0 137062 400
rect 141974 0 142030 400
rect 146942 0 146998 400
rect 152002 0 152058 400
rect 156970 0 157026 400
rect 161938 0 161994 400
rect 166906 0 166962 400
rect 171874 0 171930 400
rect 176934 0 176990 400
rect 181902 0 181958 400
rect 186870 0 186926 400
rect 191838 0 191894 400
rect 196806 0 196862 400
rect 201774 0 201830 400
rect 206834 0 206890 400
rect 211802 0 211858 400
rect 216770 0 216826 400
rect 221738 0 221794 400
rect 226706 0 226762 400
rect 231674 0 231730 400
rect 236734 0 236790 400
rect 241702 0 241758 400
rect 246670 0 246726 400
rect 251638 0 251694 400
rect 256606 0 256662 400
rect 261574 0 261630 400
rect 266634 0 266690 400
rect 271602 0 271658 400
rect 276570 0 276626 400
rect 281538 0 281594 400
rect 286506 0 286562 400
rect 291474 0 291530 400
rect 296534 0 296590 400
rect 301502 0 301558 400
rect 306470 0 306526 400
rect 311438 0 311494 400
rect 316406 0 316462 400
<< obsm2 >>
rect 296 197016 2446 197470
rect 2614 197016 7414 197470
rect 7582 197016 12382 197470
rect 12550 197016 17350 197470
rect 17518 197016 22318 197470
rect 22486 197016 27286 197470
rect 27454 197016 32346 197470
rect 32514 197016 37314 197470
rect 37482 197016 42282 197470
rect 42450 197016 47250 197470
rect 47418 197016 52218 197470
rect 52386 197016 57186 197470
rect 57354 197016 62246 197470
rect 62414 197016 67214 197470
rect 67382 197016 72182 197470
rect 72350 197016 77150 197470
rect 77318 197016 82118 197470
rect 82286 197016 87086 197470
rect 87254 197016 92146 197470
rect 92314 197016 97114 197470
rect 97282 197016 102082 197470
rect 102250 197016 107050 197470
rect 107218 197016 112018 197470
rect 112186 197016 116986 197470
rect 117154 197016 122046 197470
rect 122214 197016 127014 197470
rect 127182 197016 131982 197470
rect 132150 197016 136950 197470
rect 137118 197016 141918 197470
rect 142086 197016 146886 197470
rect 147054 197016 151946 197470
rect 152114 197016 156914 197470
rect 157082 197016 161882 197470
rect 162050 197016 166850 197470
rect 167018 197016 171818 197470
rect 171986 197016 176878 197470
rect 177046 197016 181846 197470
rect 182014 197016 186814 197470
rect 186982 197016 191782 197470
rect 191950 197016 196750 197470
rect 196918 197016 201718 197470
rect 201886 197016 206778 197470
rect 206946 197016 211746 197470
rect 211914 197016 216714 197470
rect 216882 197016 221682 197470
rect 221850 197016 226650 197470
rect 226818 197016 231618 197470
rect 231786 197016 236678 197470
rect 236846 197016 241646 197470
rect 241814 197016 246614 197470
rect 246782 197016 251582 197470
rect 251750 197016 256550 197470
rect 256718 197016 261518 197470
rect 261686 197016 266578 197470
rect 266746 197016 271546 197470
rect 271714 197016 276514 197470
rect 276682 197016 281482 197470
rect 281650 197016 286450 197470
rect 286618 197016 291418 197470
rect 291586 197016 296478 197470
rect 296646 197016 301446 197470
rect 301614 197016 306414 197470
rect 306582 197016 311382 197470
rect 311550 197016 316350 197470
rect 316518 197016 318668 197470
rect 296 456 318668 197016
rect 296 2 2446 456
rect 2614 2 7414 456
rect 7582 2 12382 456
rect 12550 2 17350 456
rect 17518 2 22318 456
rect 22486 2 27286 456
rect 27454 2 32346 456
rect 32514 2 37314 456
rect 37482 2 42282 456
rect 42450 2 47250 456
rect 47418 2 52218 456
rect 52386 2 57186 456
rect 57354 2 62246 456
rect 62414 2 67214 456
rect 67382 2 72182 456
rect 72350 2 77150 456
rect 77318 2 82118 456
rect 82286 2 87086 456
rect 87254 2 92146 456
rect 92314 2 97114 456
rect 97282 2 102082 456
rect 102250 2 107050 456
rect 107218 2 112018 456
rect 112186 2 116986 456
rect 117154 2 122046 456
rect 122214 2 127014 456
rect 127182 2 131982 456
rect 132150 2 136950 456
rect 137118 2 141918 456
rect 142086 2 146886 456
rect 147054 2 151946 456
rect 152114 2 156914 456
rect 157082 2 161882 456
rect 162050 2 166850 456
rect 167018 2 171818 456
rect 171986 2 176878 456
rect 177046 2 181846 456
rect 182014 2 186814 456
rect 186982 2 191782 456
rect 191950 2 196750 456
rect 196918 2 201718 456
rect 201886 2 206778 456
rect 206946 2 211746 456
rect 211914 2 216714 456
rect 216882 2 221682 456
rect 221850 2 226650 456
rect 226818 2 231618 456
rect 231786 2 236678 456
rect 236846 2 241646 456
rect 241814 2 246614 456
rect 246782 2 251582 456
rect 251750 2 256550 456
rect 256718 2 261518 456
rect 261686 2 266578 456
rect 266746 2 271546 456
rect 271714 2 276514 456
rect 276682 2 281482 456
rect 281650 2 286450 456
rect 286618 2 291418 456
rect 291586 2 296478 456
rect 296646 2 301446 456
rect 301614 2 306414 456
rect 306582 2 311382 456
rect 311550 2 316350 456
rect 316518 2 318668 456
<< metal3 >>
rect 318564 191904 318964 192024
rect 318564 180888 318964 181008
rect 318564 170008 318964 170128
rect 318564 158992 318964 159112
rect 318564 147976 318964 148096
rect 318564 137096 318964 137216
rect 318564 126080 318964 126200
rect 318564 115064 318964 115184
rect 318564 104184 318964 104304
rect 0 98744 400 98864
rect 318564 93168 318964 93288
rect 318564 82152 318964 82272
rect 318564 71272 318964 71392
rect 318564 60256 318964 60376
rect 318564 49240 318964 49360
rect 318564 38360 318964 38480
rect 318564 27344 318964 27464
rect 318564 16328 318964 16448
rect 318564 5448 318964 5568
<< obsm3 >>
rect 400 192104 318564 197437
rect 400 191824 318484 192104
rect 400 181088 318564 191824
rect 400 180808 318484 181088
rect 400 170208 318564 180808
rect 400 169928 318484 170208
rect 400 159192 318564 169928
rect 400 158912 318484 159192
rect 400 148176 318564 158912
rect 400 147896 318484 148176
rect 400 137296 318564 147896
rect 400 137016 318484 137296
rect 400 126280 318564 137016
rect 400 126000 318484 126280
rect 400 115264 318564 126000
rect 400 114984 318484 115264
rect 400 104384 318564 114984
rect 400 104104 318484 104384
rect 400 98944 318564 104104
rect 480 98664 318564 98944
rect 400 93368 318564 98664
rect 400 93088 318484 93368
rect 400 82352 318564 93088
rect 400 82072 318484 82352
rect 400 71472 318564 82072
rect 400 71192 318484 71472
rect 400 60456 318564 71192
rect 400 60176 318484 60456
rect 400 49440 318564 60176
rect 400 49160 318484 49440
rect 400 38560 318564 49160
rect 400 38280 318484 38560
rect 400 27544 318564 38280
rect 400 27264 318484 27544
rect 400 16528 318564 27264
rect 400 16248 318484 16528
rect 400 5648 318564 16248
rect 400 5368 318484 5648
rect 400 35 318564 5368
<< metal4 >>
rect 4738 20080 5358 177392
rect 22738 20080 23358 177392
rect 40738 20080 41358 177392
rect 58738 20080 59358 177392
rect 76738 20080 77358 177392
rect 94738 20080 95358 177392
rect 112738 20080 113358 177392
rect 130738 20080 131358 177392
rect 148738 20080 149358 177392
rect 166738 20080 167358 177392
rect 184738 20080 185358 177392
rect 202738 20080 203358 177392
rect 220738 20080 221358 177392
rect 238738 20080 239358 177392
rect 256738 20080 257358 177392
rect 274738 20080 275358 177392
rect 292738 20080 293358 177392
rect 310738 20080 311358 177392
<< obsm4 >>
rect 979 177472 313293 197437
rect 979 20000 4658 177472
rect 5438 20000 22658 177472
rect 23438 20000 40658 177472
rect 41438 20000 58658 177472
rect 59438 20000 76658 177472
rect 77438 20000 94658 177472
rect 95438 20000 112658 177472
rect 113438 20000 130658 177472
rect 131438 20000 148658 177472
rect 149438 20000 166658 177472
rect 167438 20000 184658 177472
rect 185438 20000 202658 177472
rect 203438 20000 220658 177472
rect 221438 20000 238658 177472
rect 239438 20000 256658 177472
rect 257438 20000 274658 177472
rect 275438 20000 292658 177472
rect 293438 20000 310658 177472
rect 311438 20000 313293 177472
rect 979 171 313293 20000
<< labels >>
rlabel metal3 s 318564 104184 318964 104304 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 318564 115064 318964 115184 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 318564 126080 318964 126200 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 318564 137096 318964 137216 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 318564 147976 318964 148096 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 318564 158992 318964 159112 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 318564 170008 318964 170128 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 318564 180888 318964 181008 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 318564 191904 318964 192024 6 A0[8]
port 9 nsew signal input
rlabel metal3 s 0 98744 400 98864 6 CLK
port 10 nsew signal input
rlabel metal2 s 2502 0 2558 400 6 Di0[0]
port 11 nsew signal input
rlabel metal2 s 52274 0 52330 400 6 Di0[10]
port 12 nsew signal input
rlabel metal2 s 57242 0 57298 400 6 Di0[11]
port 13 nsew signal input
rlabel metal2 s 62302 0 62358 400 6 Di0[12]
port 14 nsew signal input
rlabel metal2 s 67270 0 67326 400 6 Di0[13]
port 15 nsew signal input
rlabel metal2 s 72238 0 72294 400 6 Di0[14]
port 16 nsew signal input
rlabel metal2 s 77206 0 77262 400 6 Di0[15]
port 17 nsew signal input
rlabel metal2 s 82174 0 82230 400 6 Di0[16]
port 18 nsew signal input
rlabel metal2 s 87142 0 87198 400 6 Di0[17]
port 19 nsew signal input
rlabel metal2 s 92202 0 92258 400 6 Di0[18]
port 20 nsew signal input
rlabel metal2 s 97170 0 97226 400 6 Di0[19]
port 21 nsew signal input
rlabel metal2 s 7470 0 7526 400 6 Di0[1]
port 22 nsew signal input
rlabel metal2 s 102138 0 102194 400 6 Di0[20]
port 23 nsew signal input
rlabel metal2 s 107106 0 107162 400 6 Di0[21]
port 24 nsew signal input
rlabel metal2 s 112074 0 112130 400 6 Di0[22]
port 25 nsew signal input
rlabel metal2 s 117042 0 117098 400 6 Di0[23]
port 26 nsew signal input
rlabel metal2 s 122102 0 122158 400 6 Di0[24]
port 27 nsew signal input
rlabel metal2 s 127070 0 127126 400 6 Di0[25]
port 28 nsew signal input
rlabel metal2 s 132038 0 132094 400 6 Di0[26]
port 29 nsew signal input
rlabel metal2 s 137006 0 137062 400 6 Di0[27]
port 30 nsew signal input
rlabel metal2 s 141974 0 142030 400 6 Di0[28]
port 31 nsew signal input
rlabel metal2 s 146942 0 146998 400 6 Di0[29]
port 32 nsew signal input
rlabel metal2 s 12438 0 12494 400 6 Di0[2]
port 33 nsew signal input
rlabel metal2 s 152002 0 152058 400 6 Di0[30]
port 34 nsew signal input
rlabel metal2 s 156970 0 157026 400 6 Di0[31]
port 35 nsew signal input
rlabel metal2 s 161938 0 161994 400 6 Di0[32]
port 36 nsew signal input
rlabel metal2 s 166906 0 166962 400 6 Di0[33]
port 37 nsew signal input
rlabel metal2 s 171874 0 171930 400 6 Di0[34]
port 38 nsew signal input
rlabel metal2 s 176934 0 176990 400 6 Di0[35]
port 39 nsew signal input
rlabel metal2 s 181902 0 181958 400 6 Di0[36]
port 40 nsew signal input
rlabel metal2 s 186870 0 186926 400 6 Di0[37]
port 41 nsew signal input
rlabel metal2 s 191838 0 191894 400 6 Di0[38]
port 42 nsew signal input
rlabel metal2 s 196806 0 196862 400 6 Di0[39]
port 43 nsew signal input
rlabel metal2 s 17406 0 17462 400 6 Di0[3]
port 44 nsew signal input
rlabel metal2 s 201774 0 201830 400 6 Di0[40]
port 45 nsew signal input
rlabel metal2 s 206834 0 206890 400 6 Di0[41]
port 46 nsew signal input
rlabel metal2 s 211802 0 211858 400 6 Di0[42]
port 47 nsew signal input
rlabel metal2 s 216770 0 216826 400 6 Di0[43]
port 48 nsew signal input
rlabel metal2 s 221738 0 221794 400 6 Di0[44]
port 49 nsew signal input
rlabel metal2 s 226706 0 226762 400 6 Di0[45]
port 50 nsew signal input
rlabel metal2 s 231674 0 231730 400 6 Di0[46]
port 51 nsew signal input
rlabel metal2 s 236734 0 236790 400 6 Di0[47]
port 52 nsew signal input
rlabel metal2 s 241702 0 241758 400 6 Di0[48]
port 53 nsew signal input
rlabel metal2 s 246670 0 246726 400 6 Di0[49]
port 54 nsew signal input
rlabel metal2 s 22374 0 22430 400 6 Di0[4]
port 55 nsew signal input
rlabel metal2 s 251638 0 251694 400 6 Di0[50]
port 56 nsew signal input
rlabel metal2 s 256606 0 256662 400 6 Di0[51]
port 57 nsew signal input
rlabel metal2 s 261574 0 261630 400 6 Di0[52]
port 58 nsew signal input
rlabel metal2 s 266634 0 266690 400 6 Di0[53]
port 59 nsew signal input
rlabel metal2 s 271602 0 271658 400 6 Di0[54]
port 60 nsew signal input
rlabel metal2 s 276570 0 276626 400 6 Di0[55]
port 61 nsew signal input
rlabel metal2 s 281538 0 281594 400 6 Di0[56]
port 62 nsew signal input
rlabel metal2 s 286506 0 286562 400 6 Di0[57]
port 63 nsew signal input
rlabel metal2 s 291474 0 291530 400 6 Di0[58]
port 64 nsew signal input
rlabel metal2 s 296534 0 296590 400 6 Di0[59]
port 65 nsew signal input
rlabel metal2 s 27342 0 27398 400 6 Di0[5]
port 66 nsew signal input
rlabel metal2 s 301502 0 301558 400 6 Di0[60]
port 67 nsew signal input
rlabel metal2 s 306470 0 306526 400 6 Di0[61]
port 68 nsew signal input
rlabel metal2 s 311438 0 311494 400 6 Di0[62]
port 69 nsew signal input
rlabel metal2 s 316406 0 316462 400 6 Di0[63]
port 70 nsew signal input
rlabel metal2 s 32402 0 32458 400 6 Di0[6]
port 71 nsew signal input
rlabel metal2 s 37370 0 37426 400 6 Di0[7]
port 72 nsew signal input
rlabel metal2 s 42338 0 42394 400 6 Di0[8]
port 73 nsew signal input
rlabel metal2 s 47306 0 47362 400 6 Di0[9]
port 74 nsew signal input
rlabel metal2 s 2502 197072 2558 197472 6 Do0[0]
port 75 nsew signal output
rlabel metal2 s 52274 197072 52330 197472 6 Do0[10]
port 76 nsew signal output
rlabel metal2 s 57242 197072 57298 197472 6 Do0[11]
port 77 nsew signal output
rlabel metal2 s 62302 197072 62358 197472 6 Do0[12]
port 78 nsew signal output
rlabel metal2 s 67270 197072 67326 197472 6 Do0[13]
port 79 nsew signal output
rlabel metal2 s 72238 197072 72294 197472 6 Do0[14]
port 80 nsew signal output
rlabel metal2 s 77206 197072 77262 197472 6 Do0[15]
port 81 nsew signal output
rlabel metal2 s 82174 197072 82230 197472 6 Do0[16]
port 82 nsew signal output
rlabel metal2 s 87142 197072 87198 197472 6 Do0[17]
port 83 nsew signal output
rlabel metal2 s 92202 197072 92258 197472 6 Do0[18]
port 84 nsew signal output
rlabel metal2 s 97170 197072 97226 197472 6 Do0[19]
port 85 nsew signal output
rlabel metal2 s 7470 197072 7526 197472 6 Do0[1]
port 86 nsew signal output
rlabel metal2 s 102138 197072 102194 197472 6 Do0[20]
port 87 nsew signal output
rlabel metal2 s 107106 197072 107162 197472 6 Do0[21]
port 88 nsew signal output
rlabel metal2 s 112074 197072 112130 197472 6 Do0[22]
port 89 nsew signal output
rlabel metal2 s 117042 197072 117098 197472 6 Do0[23]
port 90 nsew signal output
rlabel metal2 s 122102 197072 122158 197472 6 Do0[24]
port 91 nsew signal output
rlabel metal2 s 127070 197072 127126 197472 6 Do0[25]
port 92 nsew signal output
rlabel metal2 s 132038 197072 132094 197472 6 Do0[26]
port 93 nsew signal output
rlabel metal2 s 137006 197072 137062 197472 6 Do0[27]
port 94 nsew signal output
rlabel metal2 s 141974 197072 142030 197472 6 Do0[28]
port 95 nsew signal output
rlabel metal2 s 146942 197072 146998 197472 6 Do0[29]
port 96 nsew signal output
rlabel metal2 s 12438 197072 12494 197472 6 Do0[2]
port 97 nsew signal output
rlabel metal2 s 152002 197072 152058 197472 6 Do0[30]
port 98 nsew signal output
rlabel metal2 s 156970 197072 157026 197472 6 Do0[31]
port 99 nsew signal output
rlabel metal2 s 161938 197072 161994 197472 6 Do0[32]
port 100 nsew signal output
rlabel metal2 s 166906 197072 166962 197472 6 Do0[33]
port 101 nsew signal output
rlabel metal2 s 171874 197072 171930 197472 6 Do0[34]
port 102 nsew signal output
rlabel metal2 s 176934 197072 176990 197472 6 Do0[35]
port 103 nsew signal output
rlabel metal2 s 181902 197072 181958 197472 6 Do0[36]
port 104 nsew signal output
rlabel metal2 s 186870 197072 186926 197472 6 Do0[37]
port 105 nsew signal output
rlabel metal2 s 191838 197072 191894 197472 6 Do0[38]
port 106 nsew signal output
rlabel metal2 s 196806 197072 196862 197472 6 Do0[39]
port 107 nsew signal output
rlabel metal2 s 17406 197072 17462 197472 6 Do0[3]
port 108 nsew signal output
rlabel metal2 s 201774 197072 201830 197472 6 Do0[40]
port 109 nsew signal output
rlabel metal2 s 206834 197072 206890 197472 6 Do0[41]
port 110 nsew signal output
rlabel metal2 s 211802 197072 211858 197472 6 Do0[42]
port 111 nsew signal output
rlabel metal2 s 216770 197072 216826 197472 6 Do0[43]
port 112 nsew signal output
rlabel metal2 s 221738 197072 221794 197472 6 Do0[44]
port 113 nsew signal output
rlabel metal2 s 226706 197072 226762 197472 6 Do0[45]
port 114 nsew signal output
rlabel metal2 s 231674 197072 231730 197472 6 Do0[46]
port 115 nsew signal output
rlabel metal2 s 236734 197072 236790 197472 6 Do0[47]
port 116 nsew signal output
rlabel metal2 s 241702 197072 241758 197472 6 Do0[48]
port 117 nsew signal output
rlabel metal2 s 246670 197072 246726 197472 6 Do0[49]
port 118 nsew signal output
rlabel metal2 s 22374 197072 22430 197472 6 Do0[4]
port 119 nsew signal output
rlabel metal2 s 251638 197072 251694 197472 6 Do0[50]
port 120 nsew signal output
rlabel metal2 s 256606 197072 256662 197472 6 Do0[51]
port 121 nsew signal output
rlabel metal2 s 261574 197072 261630 197472 6 Do0[52]
port 122 nsew signal output
rlabel metal2 s 266634 197072 266690 197472 6 Do0[53]
port 123 nsew signal output
rlabel metal2 s 271602 197072 271658 197472 6 Do0[54]
port 124 nsew signal output
rlabel metal2 s 276570 197072 276626 197472 6 Do0[55]
port 125 nsew signal output
rlabel metal2 s 281538 197072 281594 197472 6 Do0[56]
port 126 nsew signal output
rlabel metal2 s 286506 197072 286562 197472 6 Do0[57]
port 127 nsew signal output
rlabel metal2 s 291474 197072 291530 197472 6 Do0[58]
port 128 nsew signal output
rlabel metal2 s 296534 197072 296590 197472 6 Do0[59]
port 129 nsew signal output
rlabel metal2 s 27342 197072 27398 197472 6 Do0[5]
port 130 nsew signal output
rlabel metal2 s 301502 197072 301558 197472 6 Do0[60]
port 131 nsew signal output
rlabel metal2 s 306470 197072 306526 197472 6 Do0[61]
port 132 nsew signal output
rlabel metal2 s 311438 197072 311494 197472 6 Do0[62]
port 133 nsew signal output
rlabel metal2 s 316406 197072 316462 197472 6 Do0[63]
port 134 nsew signal output
rlabel metal2 s 32402 197072 32458 197472 6 Do0[6]
port 135 nsew signal output
rlabel metal2 s 37370 197072 37426 197472 6 Do0[7]
port 136 nsew signal output
rlabel metal2 s 42338 197072 42394 197472 6 Do0[8]
port 137 nsew signal output
rlabel metal2 s 47306 197072 47362 197472 6 Do0[9]
port 138 nsew signal output
rlabel metal3 s 318564 5448 318964 5568 6 EN0
port 139 nsew signal input
rlabel metal4 s 22738 20080 23358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 58738 20080 59358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 94738 20080 95358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 130738 20080 131358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 166738 20080 167358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 202738 20080 203358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 238738 20080 239358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 274738 20080 275358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 310738 20080 311358 177392 6 VGND
port 140 nsew ground input
rlabel metal4 s 4738 20080 5358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 40738 20080 41358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 76738 20080 77358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 112738 20080 113358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 148738 20080 149358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 184738 20080 185358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 220738 20080 221358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 256738 20080 257358 177392 6 VPWR
port 141 nsew power input
rlabel metal4 s 292738 20080 293358 177392 6 VPWR
port 141 nsew power input
rlabel metal3 s 318564 16328 318964 16448 6 WE0[0]
port 142 nsew signal input
rlabel metal3 s 318564 27344 318964 27464 6 WE0[1]
port 143 nsew signal input
rlabel metal3 s 318564 38360 318964 38480 6 WE0[2]
port 144 nsew signal input
rlabel metal3 s 318564 49240 318964 49360 6 WE0[3]
port 145 nsew signal input
rlabel metal3 s 318564 60256 318964 60376 6 WE0[4]
port 146 nsew signal input
rlabel metal3 s 318564 71272 318964 71392 6 WE0[5]
port 147 nsew signal input
rlabel metal3 s 318564 82152 318964 82272 6 WE0[6]
port 148 nsew signal input
rlabel metal3 s 318564 93168 318964 93288 6 WE0[7]
port 149 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 318964 197472
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 194242612
string GDS_FILE /mnt/dffram/build/512x64_DEFAULT/openlane/runs/RUN_2022.02.20_09.14.56/results/finishing/RAM512.magic.gds
string GDS_START 165654
<< end >>

