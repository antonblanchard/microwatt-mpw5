magic
tech sky130A
magscale 1 2
timestamp 1647886595
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 198 1980 110000 107760
<< metal2 >>
rect 386 109200 442 110000
rect 1214 109200 1270 110000
rect 2042 109200 2098 110000
rect 2870 109200 2926 110000
rect 3698 109200 3754 110000
rect 4618 109200 4674 110000
rect 5446 109200 5502 110000
rect 6274 109200 6330 110000
rect 7102 109200 7158 110000
rect 7930 109200 7986 110000
rect 8850 109200 8906 110000
rect 9678 109200 9734 110000
rect 10506 109200 10562 110000
rect 11334 109200 11390 110000
rect 12162 109200 12218 110000
rect 13082 109200 13138 110000
rect 13910 109200 13966 110000
rect 14738 109200 14794 110000
rect 15566 109200 15622 110000
rect 16394 109200 16450 110000
rect 17314 109200 17370 110000
rect 18142 109200 18198 110000
rect 18970 109200 19026 110000
rect 19798 109200 19854 110000
rect 20626 109200 20682 110000
rect 21546 109200 21602 110000
rect 22374 109200 22430 110000
rect 23202 109200 23258 110000
rect 24030 109200 24086 110000
rect 24858 109200 24914 110000
rect 25778 109200 25834 110000
rect 26606 109200 26662 110000
rect 27434 109200 27490 110000
rect 28262 109200 28318 110000
rect 29090 109200 29146 110000
rect 30010 109200 30066 110000
rect 30838 109200 30894 110000
rect 31666 109200 31722 110000
rect 32494 109200 32550 110000
rect 33322 109200 33378 110000
rect 34242 109200 34298 110000
rect 35070 109200 35126 110000
rect 35898 109200 35954 110000
rect 36726 109200 36782 110000
rect 37554 109200 37610 110000
rect 38474 109200 38530 110000
rect 39302 109200 39358 110000
rect 40130 109200 40186 110000
rect 40958 109200 41014 110000
rect 41786 109200 41842 110000
rect 42706 109200 42762 110000
rect 43534 109200 43590 110000
rect 44362 109200 44418 110000
rect 45190 109200 45246 110000
rect 46018 109200 46074 110000
rect 46938 109200 46994 110000
rect 47766 109200 47822 110000
rect 48594 109200 48650 110000
rect 49422 109200 49478 110000
rect 50250 109200 50306 110000
rect 51170 109200 51226 110000
rect 51998 109200 52054 110000
rect 52826 109200 52882 110000
rect 53654 109200 53710 110000
rect 54482 109200 54538 110000
rect 55402 109200 55458 110000
rect 56230 109200 56286 110000
rect 57058 109200 57114 110000
rect 57886 109200 57942 110000
rect 58714 109200 58770 110000
rect 59634 109200 59690 110000
rect 60462 109200 60518 110000
rect 61290 109200 61346 110000
rect 62118 109200 62174 110000
rect 62946 109200 63002 110000
rect 63866 109200 63922 110000
rect 64694 109200 64750 110000
rect 65522 109200 65578 110000
rect 66350 109200 66406 110000
rect 67178 109200 67234 110000
rect 68098 109200 68154 110000
rect 68926 109200 68982 110000
rect 69754 109200 69810 110000
rect 70582 109200 70638 110000
rect 71410 109200 71466 110000
rect 72330 109200 72386 110000
rect 73158 109200 73214 110000
rect 73986 109200 74042 110000
rect 74814 109200 74870 110000
rect 75642 109200 75698 110000
rect 76562 109200 76618 110000
rect 77390 109200 77446 110000
rect 78218 109200 78274 110000
rect 79046 109200 79102 110000
rect 79874 109200 79930 110000
rect 80794 109200 80850 110000
rect 81622 109200 81678 110000
rect 82450 109200 82506 110000
rect 83278 109200 83334 110000
rect 84106 109200 84162 110000
rect 85026 109200 85082 110000
rect 85854 109200 85910 110000
rect 86682 109200 86738 110000
rect 87510 109200 87566 110000
rect 88338 109200 88394 110000
rect 89258 109200 89314 110000
rect 90086 109200 90142 110000
rect 90914 109200 90970 110000
rect 91742 109200 91798 110000
rect 92570 109200 92626 110000
rect 93490 109200 93546 110000
rect 94318 109200 94374 110000
rect 95146 109200 95202 110000
rect 95974 109200 96030 110000
rect 96802 109200 96858 110000
rect 97722 109200 97778 110000
rect 98550 109200 98606 110000
rect 99378 109200 99434 110000
rect 100206 109200 100262 110000
rect 101034 109200 101090 110000
rect 101954 109200 102010 110000
rect 102782 109200 102838 110000
rect 103610 109200 103666 110000
rect 104438 109200 104494 110000
rect 105266 109200 105322 110000
rect 106186 109200 106242 110000
rect 107014 109200 107070 110000
rect 107842 109200 107898 110000
rect 108670 109200 108726 110000
rect 109498 109200 109554 110000
rect 386 0 442 800
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2962 0 3018 800
rect 3790 0 3846 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7194 0 7250 800
rect 8114 0 8170 800
rect 8942 0 8998 800
rect 9770 0 9826 800
rect 10690 0 10746 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13266 0 13322 800
rect 14094 0 14150 800
rect 14922 0 14978 800
rect 15842 0 15898 800
rect 16670 0 16726 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 19246 0 19302 800
rect 20074 0 20130 800
rect 20994 0 21050 800
rect 21822 0 21878 800
rect 22650 0 22706 800
rect 23570 0 23626 800
rect 24398 0 24454 800
rect 25226 0 25282 800
rect 26146 0 26202 800
rect 26974 0 27030 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30470 0 30526 800
rect 31298 0 31354 800
rect 32126 0 32182 800
rect 33046 0 33102 800
rect 33874 0 33930 800
rect 34702 0 34758 800
rect 35622 0 35678 800
rect 36450 0 36506 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 39026 0 39082 800
rect 39854 0 39910 800
rect 40774 0 40830 800
rect 41602 0 41658 800
rect 42430 0 42486 800
rect 43350 0 43406 800
rect 44178 0 44234 800
rect 45006 0 45062 800
rect 45926 0 45982 800
rect 46754 0 46810 800
rect 47582 0 47638 800
rect 48502 0 48558 800
rect 49330 0 49386 800
rect 50158 0 50214 800
rect 51078 0 51134 800
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53654 0 53710 800
rect 54482 0 54538 800
rect 55402 0 55458 800
rect 56230 0 56286 800
rect 57058 0 57114 800
rect 57978 0 58034 800
rect 58806 0 58862 800
rect 59634 0 59690 800
rect 60554 0 60610 800
rect 61382 0 61438 800
rect 62210 0 62266 800
rect 63130 0 63186 800
rect 63958 0 64014 800
rect 64786 0 64842 800
rect 65706 0 65762 800
rect 66534 0 66590 800
rect 67362 0 67418 800
rect 68282 0 68338 800
rect 69110 0 69166 800
rect 69938 0 69994 800
rect 70858 0 70914 800
rect 71686 0 71742 800
rect 72514 0 72570 800
rect 73434 0 73490 800
rect 74262 0 74318 800
rect 75090 0 75146 800
rect 76010 0 76066 800
rect 76838 0 76894 800
rect 77666 0 77722 800
rect 78586 0 78642 800
rect 79414 0 79470 800
rect 80242 0 80298 800
rect 81162 0 81218 800
rect 81990 0 82046 800
rect 82910 0 82966 800
rect 83738 0 83794 800
rect 84566 0 84622 800
rect 85486 0 85542 800
rect 86314 0 86370 800
rect 87142 0 87198 800
rect 88062 0 88118 800
rect 88890 0 88946 800
rect 89718 0 89774 800
rect 90638 0 90694 800
rect 91466 0 91522 800
rect 92294 0 92350 800
rect 93214 0 93270 800
rect 94042 0 94098 800
rect 94870 0 94926 800
rect 95790 0 95846 800
rect 96618 0 96674 800
rect 97446 0 97502 800
rect 98366 0 98422 800
rect 99194 0 99250 800
rect 100022 0 100078 800
rect 100942 0 100998 800
rect 101770 0 101826 800
rect 102598 0 102654 800
rect 103518 0 103574 800
rect 104346 0 104402 800
rect 105174 0 105230 800
rect 106094 0 106150 800
rect 106922 0 106978 800
rect 107750 0 107806 800
rect 108670 0 108726 800
rect 109498 0 109554 800
<< obsm2 >>
rect 202 109144 330 109585
rect 498 109144 1158 109585
rect 1326 109144 1986 109585
rect 2154 109144 2814 109585
rect 2982 109144 3642 109585
rect 3810 109144 4562 109585
rect 4730 109144 5390 109585
rect 5558 109144 6218 109585
rect 6386 109144 7046 109585
rect 7214 109144 7874 109585
rect 8042 109144 8794 109585
rect 8962 109144 9622 109585
rect 9790 109144 10450 109585
rect 10618 109144 11278 109585
rect 11446 109144 12106 109585
rect 12274 109144 13026 109585
rect 13194 109144 13854 109585
rect 14022 109144 14682 109585
rect 14850 109144 15510 109585
rect 15678 109144 16338 109585
rect 16506 109144 17258 109585
rect 17426 109144 18086 109585
rect 18254 109144 18914 109585
rect 19082 109144 19742 109585
rect 19910 109144 20570 109585
rect 20738 109144 21490 109585
rect 21658 109144 22318 109585
rect 22486 109144 23146 109585
rect 23314 109144 23974 109585
rect 24142 109144 24802 109585
rect 24970 109144 25722 109585
rect 25890 109144 26550 109585
rect 26718 109144 27378 109585
rect 27546 109144 28206 109585
rect 28374 109144 29034 109585
rect 29202 109144 29954 109585
rect 30122 109144 30782 109585
rect 30950 109144 31610 109585
rect 31778 109144 32438 109585
rect 32606 109144 33266 109585
rect 33434 109144 34186 109585
rect 34354 109144 35014 109585
rect 35182 109144 35842 109585
rect 36010 109144 36670 109585
rect 36838 109144 37498 109585
rect 37666 109144 38418 109585
rect 38586 109144 39246 109585
rect 39414 109144 40074 109585
rect 40242 109144 40902 109585
rect 41070 109144 41730 109585
rect 41898 109144 42650 109585
rect 42818 109144 43478 109585
rect 43646 109144 44306 109585
rect 44474 109144 45134 109585
rect 45302 109144 45962 109585
rect 46130 109144 46882 109585
rect 47050 109144 47710 109585
rect 47878 109144 48538 109585
rect 48706 109144 49366 109585
rect 49534 109144 50194 109585
rect 50362 109144 51114 109585
rect 51282 109144 51942 109585
rect 52110 109144 52770 109585
rect 52938 109144 53598 109585
rect 53766 109144 54426 109585
rect 54594 109144 55346 109585
rect 55514 109144 56174 109585
rect 56342 109144 57002 109585
rect 57170 109144 57830 109585
rect 57998 109144 58658 109585
rect 58826 109144 59578 109585
rect 59746 109144 60406 109585
rect 60574 109144 61234 109585
rect 61402 109144 62062 109585
rect 62230 109144 62890 109585
rect 63058 109144 63810 109585
rect 63978 109144 64638 109585
rect 64806 109144 65466 109585
rect 65634 109144 66294 109585
rect 66462 109144 67122 109585
rect 67290 109144 68042 109585
rect 68210 109144 68870 109585
rect 69038 109144 69698 109585
rect 69866 109144 70526 109585
rect 70694 109144 71354 109585
rect 71522 109144 72274 109585
rect 72442 109144 73102 109585
rect 73270 109144 73930 109585
rect 74098 109144 74758 109585
rect 74926 109144 75586 109585
rect 75754 109144 76506 109585
rect 76674 109144 77334 109585
rect 77502 109144 78162 109585
rect 78330 109144 78990 109585
rect 79158 109144 79818 109585
rect 79986 109144 80738 109585
rect 80906 109144 81566 109585
rect 81734 109144 82394 109585
rect 82562 109144 83222 109585
rect 83390 109144 84050 109585
rect 84218 109144 84970 109585
rect 85138 109144 85798 109585
rect 85966 109144 86626 109585
rect 86794 109144 87454 109585
rect 87622 109144 88282 109585
rect 88450 109144 89202 109585
rect 89370 109144 90030 109585
rect 90198 109144 90858 109585
rect 91026 109144 91686 109585
rect 91854 109144 92514 109585
rect 92682 109144 93434 109585
rect 93602 109144 94262 109585
rect 94430 109144 95090 109585
rect 95258 109144 95918 109585
rect 96086 109144 96746 109585
rect 96914 109144 97666 109585
rect 97834 109144 98494 109585
rect 98662 109144 99322 109585
rect 99490 109144 100150 109585
rect 100318 109144 100978 109585
rect 101146 109144 101898 109585
rect 102066 109144 102726 109585
rect 102894 109144 103554 109585
rect 103722 109144 104382 109585
rect 104550 109144 105210 109585
rect 105378 109144 106130 109585
rect 106298 109144 106958 109585
rect 107126 109144 107786 109585
rect 107954 109144 108614 109585
rect 108782 109144 109442 109585
rect 109610 109144 110000 109585
rect 202 856 110000 109144
rect 202 439 330 856
rect 498 439 1158 856
rect 1326 439 1986 856
rect 2154 439 2906 856
rect 3074 439 3734 856
rect 3902 439 4562 856
rect 4730 439 5482 856
rect 5650 439 6310 856
rect 6478 439 7138 856
rect 7306 439 8058 856
rect 8226 439 8886 856
rect 9054 439 9714 856
rect 9882 439 10634 856
rect 10802 439 11462 856
rect 11630 439 12290 856
rect 12458 439 13210 856
rect 13378 439 14038 856
rect 14206 439 14866 856
rect 15034 439 15786 856
rect 15954 439 16614 856
rect 16782 439 17442 856
rect 17610 439 18362 856
rect 18530 439 19190 856
rect 19358 439 20018 856
rect 20186 439 20938 856
rect 21106 439 21766 856
rect 21934 439 22594 856
rect 22762 439 23514 856
rect 23682 439 24342 856
rect 24510 439 25170 856
rect 25338 439 26090 856
rect 26258 439 26918 856
rect 27086 439 27838 856
rect 28006 439 28666 856
rect 28834 439 29494 856
rect 29662 439 30414 856
rect 30582 439 31242 856
rect 31410 439 32070 856
rect 32238 439 32990 856
rect 33158 439 33818 856
rect 33986 439 34646 856
rect 34814 439 35566 856
rect 35734 439 36394 856
rect 36562 439 37222 856
rect 37390 439 38142 856
rect 38310 439 38970 856
rect 39138 439 39798 856
rect 39966 439 40718 856
rect 40886 439 41546 856
rect 41714 439 42374 856
rect 42542 439 43294 856
rect 43462 439 44122 856
rect 44290 439 44950 856
rect 45118 439 45870 856
rect 46038 439 46698 856
rect 46866 439 47526 856
rect 47694 439 48446 856
rect 48614 439 49274 856
rect 49442 439 50102 856
rect 50270 439 51022 856
rect 51190 439 51850 856
rect 52018 439 52678 856
rect 52846 439 53598 856
rect 53766 439 54426 856
rect 54594 439 55346 856
rect 55514 439 56174 856
rect 56342 439 57002 856
rect 57170 439 57922 856
rect 58090 439 58750 856
rect 58918 439 59578 856
rect 59746 439 60498 856
rect 60666 439 61326 856
rect 61494 439 62154 856
rect 62322 439 63074 856
rect 63242 439 63902 856
rect 64070 439 64730 856
rect 64898 439 65650 856
rect 65818 439 66478 856
rect 66646 439 67306 856
rect 67474 439 68226 856
rect 68394 439 69054 856
rect 69222 439 69882 856
rect 70050 439 70802 856
rect 70970 439 71630 856
rect 71798 439 72458 856
rect 72626 439 73378 856
rect 73546 439 74206 856
rect 74374 439 75034 856
rect 75202 439 75954 856
rect 76122 439 76782 856
rect 76950 439 77610 856
rect 77778 439 78530 856
rect 78698 439 79358 856
rect 79526 439 80186 856
rect 80354 439 81106 856
rect 81274 439 81934 856
rect 82102 439 82854 856
rect 83022 439 83682 856
rect 83850 439 84510 856
rect 84678 439 85430 856
rect 85598 439 86258 856
rect 86426 439 87086 856
rect 87254 439 88006 856
rect 88174 439 88834 856
rect 89002 439 89662 856
rect 89830 439 90582 856
rect 90750 439 91410 856
rect 91578 439 92238 856
rect 92406 439 93158 856
rect 93326 439 93986 856
rect 94154 439 94814 856
rect 94982 439 95734 856
rect 95902 439 96562 856
rect 96730 439 97390 856
rect 97558 439 98310 856
rect 98478 439 99138 856
rect 99306 439 99966 856
rect 100134 439 100886 856
rect 101054 439 101714 856
rect 101882 439 102542 856
rect 102710 439 103462 856
rect 103630 439 104290 856
rect 104458 439 105118 856
rect 105286 439 106038 856
rect 106206 439 106866 856
rect 107034 439 107694 856
rect 107862 439 108614 856
rect 108782 439 109442 856
rect 109610 439 110000 856
<< metal3 >>
rect 109200 109488 110000 109608
rect 109200 108672 110000 108792
rect 109200 107856 110000 107976
rect 109200 106904 110000 107024
rect 109200 106088 110000 106208
rect 109200 105272 110000 105392
rect 109200 104320 110000 104440
rect 109200 103504 110000 103624
rect 109200 102688 110000 102808
rect 109200 101736 110000 101856
rect 109200 100920 110000 101040
rect 109200 100104 110000 100224
rect 109200 99152 110000 99272
rect 109200 98336 110000 98456
rect 109200 97520 110000 97640
rect 109200 96568 110000 96688
rect 109200 95752 110000 95872
rect 109200 94936 110000 95056
rect 109200 93984 110000 94104
rect 109200 93168 110000 93288
rect 109200 92352 110000 92472
rect 109200 91400 110000 91520
rect 109200 90584 110000 90704
rect 109200 89768 110000 89888
rect 109200 88816 110000 88936
rect 109200 88000 110000 88120
rect 109200 87184 110000 87304
rect 109200 86368 110000 86488
rect 109200 85416 110000 85536
rect 109200 84600 110000 84720
rect 109200 83784 110000 83904
rect 109200 82832 110000 82952
rect 109200 82016 110000 82136
rect 109200 81200 110000 81320
rect 109200 80248 110000 80368
rect 109200 79432 110000 79552
rect 109200 78616 110000 78736
rect 109200 77664 110000 77784
rect 109200 76848 110000 76968
rect 109200 76032 110000 76152
rect 109200 75080 110000 75200
rect 109200 74264 110000 74384
rect 109200 73448 110000 73568
rect 109200 72496 110000 72616
rect 109200 71680 110000 71800
rect 109200 70864 110000 70984
rect 109200 69912 110000 70032
rect 109200 69096 110000 69216
rect 109200 68280 110000 68400
rect 109200 67328 110000 67448
rect 109200 66512 110000 66632
rect 109200 65696 110000 65816
rect 109200 64880 110000 65000
rect 109200 63928 110000 64048
rect 109200 63112 110000 63232
rect 109200 62296 110000 62416
rect 109200 61344 110000 61464
rect 109200 60528 110000 60648
rect 109200 59712 110000 59832
rect 109200 58760 110000 58880
rect 109200 57944 110000 58064
rect 109200 57128 110000 57248
rect 109200 56176 110000 56296
rect 109200 55360 110000 55480
rect 109200 54544 110000 54664
rect 109200 53592 110000 53712
rect 109200 52776 110000 52896
rect 109200 51960 110000 52080
rect 109200 51008 110000 51128
rect 109200 50192 110000 50312
rect 109200 49376 110000 49496
rect 109200 48424 110000 48544
rect 109200 47608 110000 47728
rect 109200 46792 110000 46912
rect 109200 45840 110000 45960
rect 109200 45024 110000 45144
rect 109200 44208 110000 44328
rect 109200 43392 110000 43512
rect 109200 42440 110000 42560
rect 109200 41624 110000 41744
rect 109200 40808 110000 40928
rect 109200 39856 110000 39976
rect 109200 39040 110000 39160
rect 109200 38224 110000 38344
rect 109200 37272 110000 37392
rect 109200 36456 110000 36576
rect 109200 35640 110000 35760
rect 109200 34688 110000 34808
rect 109200 33872 110000 33992
rect 109200 33056 110000 33176
rect 109200 32104 110000 32224
rect 109200 31288 110000 31408
rect 109200 30472 110000 30592
rect 109200 29520 110000 29640
rect 109200 28704 110000 28824
rect 109200 27888 110000 28008
rect 109200 26936 110000 27056
rect 109200 26120 110000 26240
rect 109200 25304 110000 25424
rect 109200 24352 110000 24472
rect 109200 23536 110000 23656
rect 109200 22720 110000 22840
rect 109200 21904 110000 22024
rect 109200 20952 110000 21072
rect 109200 20136 110000 20256
rect 109200 19320 110000 19440
rect 109200 18368 110000 18488
rect 109200 17552 110000 17672
rect 109200 16736 110000 16856
rect 109200 15784 110000 15904
rect 109200 14968 110000 15088
rect 109200 14152 110000 14272
rect 109200 13200 110000 13320
rect 109200 12384 110000 12504
rect 109200 11568 110000 11688
rect 109200 10616 110000 10736
rect 109200 9800 110000 9920
rect 109200 8984 110000 9104
rect 109200 8032 110000 8152
rect 109200 7216 110000 7336
rect 109200 6400 110000 6520
rect 109200 5448 110000 5568
rect 109200 4632 110000 4752
rect 109200 3816 110000 3936
rect 109200 2864 110000 2984
rect 109200 2048 110000 2168
rect 109200 1232 110000 1352
rect 109200 416 110000 536
<< obsm3 >>
rect 197 109408 109120 109581
rect 197 108872 109970 109408
rect 197 108592 109120 108872
rect 197 108056 109970 108592
rect 197 107776 109120 108056
rect 197 107104 109970 107776
rect 197 106824 109120 107104
rect 197 106288 109970 106824
rect 197 106008 109120 106288
rect 197 105472 109970 106008
rect 197 105192 109120 105472
rect 197 104520 109970 105192
rect 197 104240 109120 104520
rect 197 103704 109970 104240
rect 197 103424 109120 103704
rect 197 102888 109970 103424
rect 197 102608 109120 102888
rect 197 101936 109970 102608
rect 197 101656 109120 101936
rect 197 101120 109970 101656
rect 197 100840 109120 101120
rect 197 100304 109970 100840
rect 197 100024 109120 100304
rect 197 99352 109970 100024
rect 197 99072 109120 99352
rect 197 98536 109970 99072
rect 197 98256 109120 98536
rect 197 97720 109970 98256
rect 197 97440 109120 97720
rect 197 96768 109970 97440
rect 197 96488 109120 96768
rect 197 95952 109970 96488
rect 197 95672 109120 95952
rect 197 95136 109970 95672
rect 197 94856 109120 95136
rect 197 94184 109970 94856
rect 197 93904 109120 94184
rect 197 93368 109970 93904
rect 197 93088 109120 93368
rect 197 92552 109970 93088
rect 197 92272 109120 92552
rect 197 91600 109970 92272
rect 197 91320 109120 91600
rect 197 90784 109970 91320
rect 197 90504 109120 90784
rect 197 89968 109970 90504
rect 197 89688 109120 89968
rect 197 89016 109970 89688
rect 197 88736 109120 89016
rect 197 88200 109970 88736
rect 197 87920 109120 88200
rect 197 87384 109970 87920
rect 197 87104 109120 87384
rect 197 86568 109970 87104
rect 197 86288 109120 86568
rect 197 85616 109970 86288
rect 197 85336 109120 85616
rect 197 84800 109970 85336
rect 197 84520 109120 84800
rect 197 83984 109970 84520
rect 197 83704 109120 83984
rect 197 83032 109970 83704
rect 197 82752 109120 83032
rect 197 82216 109970 82752
rect 197 81936 109120 82216
rect 197 81400 109970 81936
rect 197 81120 109120 81400
rect 197 80448 109970 81120
rect 197 80168 109120 80448
rect 197 79632 109970 80168
rect 197 79352 109120 79632
rect 197 78816 109970 79352
rect 197 78536 109120 78816
rect 197 77864 109970 78536
rect 197 77584 109120 77864
rect 197 77048 109970 77584
rect 197 76768 109120 77048
rect 197 76232 109970 76768
rect 197 75952 109120 76232
rect 197 75280 109970 75952
rect 197 75000 109120 75280
rect 197 74464 109970 75000
rect 197 74184 109120 74464
rect 197 73648 109970 74184
rect 197 73368 109120 73648
rect 197 72696 109970 73368
rect 197 72416 109120 72696
rect 197 71880 109970 72416
rect 197 71600 109120 71880
rect 197 71064 109970 71600
rect 197 70784 109120 71064
rect 197 70112 109970 70784
rect 197 69832 109120 70112
rect 197 69296 109970 69832
rect 197 69016 109120 69296
rect 197 68480 109970 69016
rect 197 68200 109120 68480
rect 197 67528 109970 68200
rect 197 67248 109120 67528
rect 197 66712 109970 67248
rect 197 66432 109120 66712
rect 197 65896 109970 66432
rect 197 65616 109120 65896
rect 197 65080 109970 65616
rect 197 64800 109120 65080
rect 197 64128 109970 64800
rect 197 63848 109120 64128
rect 197 63312 109970 63848
rect 197 63032 109120 63312
rect 197 62496 109970 63032
rect 197 62216 109120 62496
rect 197 61544 109970 62216
rect 197 61264 109120 61544
rect 197 60728 109970 61264
rect 197 60448 109120 60728
rect 197 59912 109970 60448
rect 197 59632 109120 59912
rect 197 58960 109970 59632
rect 197 58680 109120 58960
rect 197 58144 109970 58680
rect 197 57864 109120 58144
rect 197 57328 109970 57864
rect 197 57048 109120 57328
rect 197 56376 109970 57048
rect 197 56096 109120 56376
rect 197 55560 109970 56096
rect 197 55280 109120 55560
rect 197 54744 109970 55280
rect 197 54464 109120 54744
rect 197 53792 109970 54464
rect 197 53512 109120 53792
rect 197 52976 109970 53512
rect 197 52696 109120 52976
rect 197 52160 109970 52696
rect 197 51880 109120 52160
rect 197 51208 109970 51880
rect 197 50928 109120 51208
rect 197 50392 109970 50928
rect 197 50112 109120 50392
rect 197 49576 109970 50112
rect 197 49296 109120 49576
rect 197 48624 109970 49296
rect 197 48344 109120 48624
rect 197 47808 109970 48344
rect 197 47528 109120 47808
rect 197 46992 109970 47528
rect 197 46712 109120 46992
rect 197 46040 109970 46712
rect 197 45760 109120 46040
rect 197 45224 109970 45760
rect 197 44944 109120 45224
rect 197 44408 109970 44944
rect 197 44128 109120 44408
rect 197 43592 109970 44128
rect 197 43312 109120 43592
rect 197 42640 109970 43312
rect 197 42360 109120 42640
rect 197 41824 109970 42360
rect 197 41544 109120 41824
rect 197 41008 109970 41544
rect 197 40728 109120 41008
rect 197 40056 109970 40728
rect 197 39776 109120 40056
rect 197 39240 109970 39776
rect 197 38960 109120 39240
rect 197 38424 109970 38960
rect 197 38144 109120 38424
rect 197 37472 109970 38144
rect 197 37192 109120 37472
rect 197 36656 109970 37192
rect 197 36376 109120 36656
rect 197 35840 109970 36376
rect 197 35560 109120 35840
rect 197 34888 109970 35560
rect 197 34608 109120 34888
rect 197 34072 109970 34608
rect 197 33792 109120 34072
rect 197 33256 109970 33792
rect 197 32976 109120 33256
rect 197 32304 109970 32976
rect 197 32024 109120 32304
rect 197 31488 109970 32024
rect 197 31208 109120 31488
rect 197 30672 109970 31208
rect 197 30392 109120 30672
rect 197 29720 109970 30392
rect 197 29440 109120 29720
rect 197 28904 109970 29440
rect 197 28624 109120 28904
rect 197 28088 109970 28624
rect 197 27808 109120 28088
rect 197 27136 109970 27808
rect 197 26856 109120 27136
rect 197 26320 109970 26856
rect 197 26040 109120 26320
rect 197 25504 109970 26040
rect 197 25224 109120 25504
rect 197 24552 109970 25224
rect 197 24272 109120 24552
rect 197 23736 109970 24272
rect 197 23456 109120 23736
rect 197 22920 109970 23456
rect 197 22640 109120 22920
rect 197 22104 109970 22640
rect 197 21824 109120 22104
rect 197 21152 109970 21824
rect 197 20872 109120 21152
rect 197 20336 109970 20872
rect 197 20056 109120 20336
rect 197 19520 109970 20056
rect 197 19240 109120 19520
rect 197 18568 109970 19240
rect 197 18288 109120 18568
rect 197 17752 109970 18288
rect 197 17472 109120 17752
rect 197 16936 109970 17472
rect 197 16656 109120 16936
rect 197 15984 109970 16656
rect 197 15704 109120 15984
rect 197 15168 109970 15704
rect 197 14888 109120 15168
rect 197 14352 109970 14888
rect 197 14072 109120 14352
rect 197 13400 109970 14072
rect 197 13120 109120 13400
rect 197 12584 109970 13120
rect 197 12304 109120 12584
rect 197 11768 109970 12304
rect 197 11488 109120 11768
rect 197 10816 109970 11488
rect 197 10536 109120 10816
rect 197 10000 109970 10536
rect 197 9720 109120 10000
rect 197 9184 109970 9720
rect 197 8904 109120 9184
rect 197 8232 109970 8904
rect 197 7952 109120 8232
rect 197 7416 109970 7952
rect 197 7136 109120 7416
rect 197 6600 109970 7136
rect 197 6320 109120 6600
rect 197 5648 109970 6320
rect 197 5368 109120 5648
rect 197 4832 109970 5368
rect 197 4552 109120 4832
rect 197 4016 109970 4552
rect 197 3736 109120 4016
rect 197 3064 109970 3736
rect 197 2784 109120 3064
rect 197 2248 109970 2784
rect 197 1968 109120 2248
rect 197 1432 109970 1968
rect 197 1152 109120 1432
rect 197 616 109970 1152
rect 197 443 109120 616
<< metal4 >>
rect 1794 2128 2414 107760
rect 19794 2128 20414 107760
rect 37794 2128 38414 107760
rect 55794 2128 56414 107760
rect 73794 2128 74414 107760
rect 91794 2128 92414 107760
<< obsm4 >>
rect 427 2048 1714 107541
rect 2494 2048 19714 107541
rect 20494 2048 37714 107541
rect 38494 2048 55714 107541
rect 56494 2048 73714 107541
rect 74494 2048 91714 107541
rect 92494 2048 108133 107541
rect 427 1667 108133 2048
<< labels >>
rlabel metal4 s 19794 2128 20414 107760 6 VGND
port 1 nsew ground input
rlabel metal4 s 55794 2128 56414 107760 6 VGND
port 1 nsew ground input
rlabel metal4 s 91794 2128 92414 107760 6 VGND
port 1 nsew ground input
rlabel metal4 s 1794 2128 2414 107760 6 VPWR
port 2 nsew power input
rlabel metal4 s 37794 2128 38414 107760 6 VPWR
port 2 nsew power input
rlabel metal4 s 73794 2128 74414 107760 6 VPWR
port 2 nsew power input
rlabel metal3 s 109200 416 110000 536 6 a[0]
port 3 nsew signal input
rlabel metal3 s 109200 8984 110000 9104 6 a[10]
port 4 nsew signal input
rlabel metal3 s 109200 9800 110000 9920 6 a[11]
port 5 nsew signal input
rlabel metal3 s 109200 10616 110000 10736 6 a[12]
port 6 nsew signal input
rlabel metal3 s 109200 11568 110000 11688 6 a[13]
port 7 nsew signal input
rlabel metal3 s 109200 12384 110000 12504 6 a[14]
port 8 nsew signal input
rlabel metal3 s 109200 13200 110000 13320 6 a[15]
port 9 nsew signal input
rlabel metal3 s 109200 14152 110000 14272 6 a[16]
port 10 nsew signal input
rlabel metal3 s 109200 14968 110000 15088 6 a[17]
port 11 nsew signal input
rlabel metal3 s 109200 15784 110000 15904 6 a[18]
port 12 nsew signal input
rlabel metal3 s 109200 16736 110000 16856 6 a[19]
port 13 nsew signal input
rlabel metal3 s 109200 1232 110000 1352 6 a[1]
port 14 nsew signal input
rlabel metal3 s 109200 17552 110000 17672 6 a[20]
port 15 nsew signal input
rlabel metal3 s 109200 18368 110000 18488 6 a[21]
port 16 nsew signal input
rlabel metal3 s 109200 19320 110000 19440 6 a[22]
port 17 nsew signal input
rlabel metal3 s 109200 20136 110000 20256 6 a[23]
port 18 nsew signal input
rlabel metal3 s 109200 20952 110000 21072 6 a[24]
port 19 nsew signal input
rlabel metal3 s 109200 21904 110000 22024 6 a[25]
port 20 nsew signal input
rlabel metal3 s 109200 22720 110000 22840 6 a[26]
port 21 nsew signal input
rlabel metal3 s 109200 23536 110000 23656 6 a[27]
port 22 nsew signal input
rlabel metal3 s 109200 24352 110000 24472 6 a[28]
port 23 nsew signal input
rlabel metal3 s 109200 25304 110000 25424 6 a[29]
port 24 nsew signal input
rlabel metal3 s 109200 2048 110000 2168 6 a[2]
port 25 nsew signal input
rlabel metal3 s 109200 26120 110000 26240 6 a[30]
port 26 nsew signal input
rlabel metal3 s 109200 26936 110000 27056 6 a[31]
port 27 nsew signal input
rlabel metal3 s 109200 27888 110000 28008 6 a[32]
port 28 nsew signal input
rlabel metal3 s 109200 28704 110000 28824 6 a[33]
port 29 nsew signal input
rlabel metal3 s 109200 29520 110000 29640 6 a[34]
port 30 nsew signal input
rlabel metal3 s 109200 30472 110000 30592 6 a[35]
port 31 nsew signal input
rlabel metal3 s 109200 31288 110000 31408 6 a[36]
port 32 nsew signal input
rlabel metal3 s 109200 32104 110000 32224 6 a[37]
port 33 nsew signal input
rlabel metal3 s 109200 33056 110000 33176 6 a[38]
port 34 nsew signal input
rlabel metal3 s 109200 33872 110000 33992 6 a[39]
port 35 nsew signal input
rlabel metal3 s 109200 2864 110000 2984 6 a[3]
port 36 nsew signal input
rlabel metal3 s 109200 34688 110000 34808 6 a[40]
port 37 nsew signal input
rlabel metal3 s 109200 35640 110000 35760 6 a[41]
port 38 nsew signal input
rlabel metal3 s 109200 36456 110000 36576 6 a[42]
port 39 nsew signal input
rlabel metal3 s 109200 37272 110000 37392 6 a[43]
port 40 nsew signal input
rlabel metal3 s 109200 38224 110000 38344 6 a[44]
port 41 nsew signal input
rlabel metal3 s 109200 39040 110000 39160 6 a[45]
port 42 nsew signal input
rlabel metal3 s 109200 39856 110000 39976 6 a[46]
port 43 nsew signal input
rlabel metal3 s 109200 40808 110000 40928 6 a[47]
port 44 nsew signal input
rlabel metal3 s 109200 41624 110000 41744 6 a[48]
port 45 nsew signal input
rlabel metal3 s 109200 42440 110000 42560 6 a[49]
port 46 nsew signal input
rlabel metal3 s 109200 3816 110000 3936 6 a[4]
port 47 nsew signal input
rlabel metal3 s 109200 43392 110000 43512 6 a[50]
port 48 nsew signal input
rlabel metal3 s 109200 44208 110000 44328 6 a[51]
port 49 nsew signal input
rlabel metal3 s 109200 45024 110000 45144 6 a[52]
port 50 nsew signal input
rlabel metal3 s 109200 45840 110000 45960 6 a[53]
port 51 nsew signal input
rlabel metal3 s 109200 46792 110000 46912 6 a[54]
port 52 nsew signal input
rlabel metal3 s 109200 47608 110000 47728 6 a[55]
port 53 nsew signal input
rlabel metal3 s 109200 48424 110000 48544 6 a[56]
port 54 nsew signal input
rlabel metal3 s 109200 49376 110000 49496 6 a[57]
port 55 nsew signal input
rlabel metal3 s 109200 50192 110000 50312 6 a[58]
port 56 nsew signal input
rlabel metal3 s 109200 51008 110000 51128 6 a[59]
port 57 nsew signal input
rlabel metal3 s 109200 4632 110000 4752 6 a[5]
port 58 nsew signal input
rlabel metal3 s 109200 51960 110000 52080 6 a[60]
port 59 nsew signal input
rlabel metal3 s 109200 52776 110000 52896 6 a[61]
port 60 nsew signal input
rlabel metal3 s 109200 53592 110000 53712 6 a[62]
port 61 nsew signal input
rlabel metal3 s 109200 54544 110000 54664 6 a[63]
port 62 nsew signal input
rlabel metal3 s 109200 5448 110000 5568 6 a[6]
port 63 nsew signal input
rlabel metal3 s 109200 6400 110000 6520 6 a[7]
port 64 nsew signal input
rlabel metal3 s 109200 7216 110000 7336 6 a[8]
port 65 nsew signal input
rlabel metal3 s 109200 8032 110000 8152 6 a[9]
port 66 nsew signal input
rlabel metal3 s 109200 55360 110000 55480 6 b[0]
port 67 nsew signal input
rlabel metal3 s 109200 63928 110000 64048 6 b[10]
port 68 nsew signal input
rlabel metal3 s 109200 64880 110000 65000 6 b[11]
port 69 nsew signal input
rlabel metal3 s 109200 65696 110000 65816 6 b[12]
port 70 nsew signal input
rlabel metal3 s 109200 66512 110000 66632 6 b[13]
port 71 nsew signal input
rlabel metal3 s 109200 67328 110000 67448 6 b[14]
port 72 nsew signal input
rlabel metal3 s 109200 68280 110000 68400 6 b[15]
port 73 nsew signal input
rlabel metal3 s 109200 69096 110000 69216 6 b[16]
port 74 nsew signal input
rlabel metal3 s 109200 69912 110000 70032 6 b[17]
port 75 nsew signal input
rlabel metal3 s 109200 70864 110000 70984 6 b[18]
port 76 nsew signal input
rlabel metal3 s 109200 71680 110000 71800 6 b[19]
port 77 nsew signal input
rlabel metal3 s 109200 56176 110000 56296 6 b[1]
port 78 nsew signal input
rlabel metal3 s 109200 72496 110000 72616 6 b[20]
port 79 nsew signal input
rlabel metal3 s 109200 73448 110000 73568 6 b[21]
port 80 nsew signal input
rlabel metal3 s 109200 74264 110000 74384 6 b[22]
port 81 nsew signal input
rlabel metal3 s 109200 75080 110000 75200 6 b[23]
port 82 nsew signal input
rlabel metal3 s 109200 76032 110000 76152 6 b[24]
port 83 nsew signal input
rlabel metal3 s 109200 76848 110000 76968 6 b[25]
port 84 nsew signal input
rlabel metal3 s 109200 77664 110000 77784 6 b[26]
port 85 nsew signal input
rlabel metal3 s 109200 78616 110000 78736 6 b[27]
port 86 nsew signal input
rlabel metal3 s 109200 79432 110000 79552 6 b[28]
port 87 nsew signal input
rlabel metal3 s 109200 80248 110000 80368 6 b[29]
port 88 nsew signal input
rlabel metal3 s 109200 57128 110000 57248 6 b[2]
port 89 nsew signal input
rlabel metal3 s 109200 81200 110000 81320 6 b[30]
port 90 nsew signal input
rlabel metal3 s 109200 82016 110000 82136 6 b[31]
port 91 nsew signal input
rlabel metal3 s 109200 82832 110000 82952 6 b[32]
port 92 nsew signal input
rlabel metal3 s 109200 83784 110000 83904 6 b[33]
port 93 nsew signal input
rlabel metal3 s 109200 84600 110000 84720 6 b[34]
port 94 nsew signal input
rlabel metal3 s 109200 85416 110000 85536 6 b[35]
port 95 nsew signal input
rlabel metal3 s 109200 86368 110000 86488 6 b[36]
port 96 nsew signal input
rlabel metal3 s 109200 87184 110000 87304 6 b[37]
port 97 nsew signal input
rlabel metal3 s 109200 88000 110000 88120 6 b[38]
port 98 nsew signal input
rlabel metal3 s 109200 88816 110000 88936 6 b[39]
port 99 nsew signal input
rlabel metal3 s 109200 57944 110000 58064 6 b[3]
port 100 nsew signal input
rlabel metal3 s 109200 89768 110000 89888 6 b[40]
port 101 nsew signal input
rlabel metal3 s 109200 90584 110000 90704 6 b[41]
port 102 nsew signal input
rlabel metal3 s 109200 91400 110000 91520 6 b[42]
port 103 nsew signal input
rlabel metal3 s 109200 92352 110000 92472 6 b[43]
port 104 nsew signal input
rlabel metal3 s 109200 93168 110000 93288 6 b[44]
port 105 nsew signal input
rlabel metal3 s 109200 93984 110000 94104 6 b[45]
port 106 nsew signal input
rlabel metal3 s 109200 94936 110000 95056 6 b[46]
port 107 nsew signal input
rlabel metal3 s 109200 95752 110000 95872 6 b[47]
port 108 nsew signal input
rlabel metal3 s 109200 96568 110000 96688 6 b[48]
port 109 nsew signal input
rlabel metal3 s 109200 97520 110000 97640 6 b[49]
port 110 nsew signal input
rlabel metal3 s 109200 58760 110000 58880 6 b[4]
port 111 nsew signal input
rlabel metal3 s 109200 98336 110000 98456 6 b[50]
port 112 nsew signal input
rlabel metal3 s 109200 99152 110000 99272 6 b[51]
port 113 nsew signal input
rlabel metal3 s 109200 100104 110000 100224 6 b[52]
port 114 nsew signal input
rlabel metal3 s 109200 100920 110000 101040 6 b[53]
port 115 nsew signal input
rlabel metal3 s 109200 101736 110000 101856 6 b[54]
port 116 nsew signal input
rlabel metal3 s 109200 102688 110000 102808 6 b[55]
port 117 nsew signal input
rlabel metal3 s 109200 103504 110000 103624 6 b[56]
port 118 nsew signal input
rlabel metal3 s 109200 104320 110000 104440 6 b[57]
port 119 nsew signal input
rlabel metal3 s 109200 105272 110000 105392 6 b[58]
port 120 nsew signal input
rlabel metal3 s 109200 106088 110000 106208 6 b[59]
port 121 nsew signal input
rlabel metal3 s 109200 59712 110000 59832 6 b[5]
port 122 nsew signal input
rlabel metal3 s 109200 106904 110000 107024 6 b[60]
port 123 nsew signal input
rlabel metal3 s 109200 107856 110000 107976 6 b[61]
port 124 nsew signal input
rlabel metal3 s 109200 108672 110000 108792 6 b[62]
port 125 nsew signal input
rlabel metal3 s 109200 109488 110000 109608 6 b[63]
port 126 nsew signal input
rlabel metal3 s 109200 60528 110000 60648 6 b[6]
port 127 nsew signal input
rlabel metal3 s 109200 61344 110000 61464 6 b[7]
port 128 nsew signal input
rlabel metal3 s 109200 62296 110000 62416 6 b[8]
port 129 nsew signal input
rlabel metal3 s 109200 63112 110000 63232 6 b[9]
port 130 nsew signal input
rlabel metal2 s 386 0 442 800 6 c[0]
port 131 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 c[100]
port 132 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 c[101]
port 133 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 c[102]
port 134 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 c[103]
port 135 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 c[104]
port 136 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 c[105]
port 137 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 c[106]
port 138 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 c[107]
port 139 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 c[108]
port 140 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 c[109]
port 141 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 c[10]
port 142 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 c[110]
port 143 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 c[111]
port 144 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 c[112]
port 145 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 c[113]
port 146 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 c[114]
port 147 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 c[115]
port 148 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 c[116]
port 149 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 c[117]
port 150 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 c[118]
port 151 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 c[119]
port 152 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 c[11]
port 153 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 c[120]
port 154 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 c[121]
port 155 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 c[122]
port 156 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 c[123]
port 157 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 c[124]
port 158 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 c[125]
port 159 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 c[126]
port 160 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 c[127]
port 161 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 c[12]
port 162 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 c[13]
port 163 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 c[14]
port 164 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 c[15]
port 165 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 c[16]
port 166 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 c[17]
port 167 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 c[18]
port 168 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 c[19]
port 169 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 c[1]
port 170 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 c[20]
port 171 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 c[21]
port 172 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 c[22]
port 173 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 c[23]
port 174 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 c[24]
port 175 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 c[25]
port 176 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 c[26]
port 177 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 c[27]
port 178 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 c[28]
port 179 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 c[29]
port 180 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 c[2]
port 181 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 c[30]
port 182 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 c[31]
port 183 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 c[32]
port 184 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 c[33]
port 185 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 c[34]
port 186 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 c[35]
port 187 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 c[36]
port 188 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 c[37]
port 189 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 c[38]
port 190 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 c[39]
port 191 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 c[3]
port 192 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 c[40]
port 193 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 c[41]
port 194 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 c[42]
port 195 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 c[43]
port 196 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 c[44]
port 197 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 c[45]
port 198 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 c[46]
port 199 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 c[47]
port 200 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 c[48]
port 201 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 c[49]
port 202 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 c[4]
port 203 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 c[50]
port 204 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 c[51]
port 205 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 c[52]
port 206 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 c[53]
port 207 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 c[54]
port 208 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 c[55]
port 209 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 c[56]
port 210 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 c[57]
port 211 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 c[58]
port 212 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 c[59]
port 213 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 c[5]
port 214 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 c[60]
port 215 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 c[61]
port 216 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 c[62]
port 217 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 c[63]
port 218 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 c[64]
port 219 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 c[65]
port 220 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 c[66]
port 221 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 c[67]
port 222 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 c[68]
port 223 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 c[69]
port 224 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 c[6]
port 225 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 c[70]
port 226 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 c[71]
port 227 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 c[72]
port 228 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 c[73]
port 229 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 c[74]
port 230 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 c[75]
port 231 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 c[76]
port 232 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 c[77]
port 233 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 c[78]
port 234 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 c[79]
port 235 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 c[7]
port 236 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 c[80]
port 237 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 c[81]
port 238 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 c[82]
port 239 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 c[83]
port 240 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 c[84]
port 241 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 c[85]
port 242 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 c[86]
port 243 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 c[87]
port 244 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 c[88]
port 245 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 c[89]
port 246 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 c[8]
port 247 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 c[90]
port 248 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 c[91]
port 249 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 c[92]
port 250 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 c[93]
port 251 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 c[94]
port 252 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 c[95]
port 253 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 c[96]
port 254 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 c[97]
port 255 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 c[98]
port 256 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 c[99]
port 257 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 c[9]
port 258 nsew signal input
rlabel metal2 s 109498 109200 109554 110000 6 clk
port 259 nsew signal input
rlabel metal2 s 386 109200 442 110000 6 o[0]
port 260 nsew signal output
rlabel metal2 s 85026 109200 85082 110000 6 o[100]
port 261 nsew signal output
rlabel metal2 s 85854 109200 85910 110000 6 o[101]
port 262 nsew signal output
rlabel metal2 s 86682 109200 86738 110000 6 o[102]
port 263 nsew signal output
rlabel metal2 s 87510 109200 87566 110000 6 o[103]
port 264 nsew signal output
rlabel metal2 s 88338 109200 88394 110000 6 o[104]
port 265 nsew signal output
rlabel metal2 s 89258 109200 89314 110000 6 o[105]
port 266 nsew signal output
rlabel metal2 s 90086 109200 90142 110000 6 o[106]
port 267 nsew signal output
rlabel metal2 s 90914 109200 90970 110000 6 o[107]
port 268 nsew signal output
rlabel metal2 s 91742 109200 91798 110000 6 o[108]
port 269 nsew signal output
rlabel metal2 s 92570 109200 92626 110000 6 o[109]
port 270 nsew signal output
rlabel metal2 s 8850 109200 8906 110000 6 o[10]
port 271 nsew signal output
rlabel metal2 s 93490 109200 93546 110000 6 o[110]
port 272 nsew signal output
rlabel metal2 s 94318 109200 94374 110000 6 o[111]
port 273 nsew signal output
rlabel metal2 s 95146 109200 95202 110000 6 o[112]
port 274 nsew signal output
rlabel metal2 s 95974 109200 96030 110000 6 o[113]
port 275 nsew signal output
rlabel metal2 s 96802 109200 96858 110000 6 o[114]
port 276 nsew signal output
rlabel metal2 s 97722 109200 97778 110000 6 o[115]
port 277 nsew signal output
rlabel metal2 s 98550 109200 98606 110000 6 o[116]
port 278 nsew signal output
rlabel metal2 s 99378 109200 99434 110000 6 o[117]
port 279 nsew signal output
rlabel metal2 s 100206 109200 100262 110000 6 o[118]
port 280 nsew signal output
rlabel metal2 s 101034 109200 101090 110000 6 o[119]
port 281 nsew signal output
rlabel metal2 s 9678 109200 9734 110000 6 o[11]
port 282 nsew signal output
rlabel metal2 s 101954 109200 102010 110000 6 o[120]
port 283 nsew signal output
rlabel metal2 s 102782 109200 102838 110000 6 o[121]
port 284 nsew signal output
rlabel metal2 s 103610 109200 103666 110000 6 o[122]
port 285 nsew signal output
rlabel metal2 s 104438 109200 104494 110000 6 o[123]
port 286 nsew signal output
rlabel metal2 s 105266 109200 105322 110000 6 o[124]
port 287 nsew signal output
rlabel metal2 s 106186 109200 106242 110000 6 o[125]
port 288 nsew signal output
rlabel metal2 s 107014 109200 107070 110000 6 o[126]
port 289 nsew signal output
rlabel metal2 s 107842 109200 107898 110000 6 o[127]
port 290 nsew signal output
rlabel metal2 s 10506 109200 10562 110000 6 o[12]
port 291 nsew signal output
rlabel metal2 s 11334 109200 11390 110000 6 o[13]
port 292 nsew signal output
rlabel metal2 s 12162 109200 12218 110000 6 o[14]
port 293 nsew signal output
rlabel metal2 s 13082 109200 13138 110000 6 o[15]
port 294 nsew signal output
rlabel metal2 s 13910 109200 13966 110000 6 o[16]
port 295 nsew signal output
rlabel metal2 s 14738 109200 14794 110000 6 o[17]
port 296 nsew signal output
rlabel metal2 s 15566 109200 15622 110000 6 o[18]
port 297 nsew signal output
rlabel metal2 s 16394 109200 16450 110000 6 o[19]
port 298 nsew signal output
rlabel metal2 s 1214 109200 1270 110000 6 o[1]
port 299 nsew signal output
rlabel metal2 s 17314 109200 17370 110000 6 o[20]
port 300 nsew signal output
rlabel metal2 s 18142 109200 18198 110000 6 o[21]
port 301 nsew signal output
rlabel metal2 s 18970 109200 19026 110000 6 o[22]
port 302 nsew signal output
rlabel metal2 s 19798 109200 19854 110000 6 o[23]
port 303 nsew signal output
rlabel metal2 s 20626 109200 20682 110000 6 o[24]
port 304 nsew signal output
rlabel metal2 s 21546 109200 21602 110000 6 o[25]
port 305 nsew signal output
rlabel metal2 s 22374 109200 22430 110000 6 o[26]
port 306 nsew signal output
rlabel metal2 s 23202 109200 23258 110000 6 o[27]
port 307 nsew signal output
rlabel metal2 s 24030 109200 24086 110000 6 o[28]
port 308 nsew signal output
rlabel metal2 s 24858 109200 24914 110000 6 o[29]
port 309 nsew signal output
rlabel metal2 s 2042 109200 2098 110000 6 o[2]
port 310 nsew signal output
rlabel metal2 s 25778 109200 25834 110000 6 o[30]
port 311 nsew signal output
rlabel metal2 s 26606 109200 26662 110000 6 o[31]
port 312 nsew signal output
rlabel metal2 s 27434 109200 27490 110000 6 o[32]
port 313 nsew signal output
rlabel metal2 s 28262 109200 28318 110000 6 o[33]
port 314 nsew signal output
rlabel metal2 s 29090 109200 29146 110000 6 o[34]
port 315 nsew signal output
rlabel metal2 s 30010 109200 30066 110000 6 o[35]
port 316 nsew signal output
rlabel metal2 s 30838 109200 30894 110000 6 o[36]
port 317 nsew signal output
rlabel metal2 s 31666 109200 31722 110000 6 o[37]
port 318 nsew signal output
rlabel metal2 s 32494 109200 32550 110000 6 o[38]
port 319 nsew signal output
rlabel metal2 s 33322 109200 33378 110000 6 o[39]
port 320 nsew signal output
rlabel metal2 s 2870 109200 2926 110000 6 o[3]
port 321 nsew signal output
rlabel metal2 s 34242 109200 34298 110000 6 o[40]
port 322 nsew signal output
rlabel metal2 s 35070 109200 35126 110000 6 o[41]
port 323 nsew signal output
rlabel metal2 s 35898 109200 35954 110000 6 o[42]
port 324 nsew signal output
rlabel metal2 s 36726 109200 36782 110000 6 o[43]
port 325 nsew signal output
rlabel metal2 s 37554 109200 37610 110000 6 o[44]
port 326 nsew signal output
rlabel metal2 s 38474 109200 38530 110000 6 o[45]
port 327 nsew signal output
rlabel metal2 s 39302 109200 39358 110000 6 o[46]
port 328 nsew signal output
rlabel metal2 s 40130 109200 40186 110000 6 o[47]
port 329 nsew signal output
rlabel metal2 s 40958 109200 41014 110000 6 o[48]
port 330 nsew signal output
rlabel metal2 s 41786 109200 41842 110000 6 o[49]
port 331 nsew signal output
rlabel metal2 s 3698 109200 3754 110000 6 o[4]
port 332 nsew signal output
rlabel metal2 s 42706 109200 42762 110000 6 o[50]
port 333 nsew signal output
rlabel metal2 s 43534 109200 43590 110000 6 o[51]
port 334 nsew signal output
rlabel metal2 s 44362 109200 44418 110000 6 o[52]
port 335 nsew signal output
rlabel metal2 s 45190 109200 45246 110000 6 o[53]
port 336 nsew signal output
rlabel metal2 s 46018 109200 46074 110000 6 o[54]
port 337 nsew signal output
rlabel metal2 s 46938 109200 46994 110000 6 o[55]
port 338 nsew signal output
rlabel metal2 s 47766 109200 47822 110000 6 o[56]
port 339 nsew signal output
rlabel metal2 s 48594 109200 48650 110000 6 o[57]
port 340 nsew signal output
rlabel metal2 s 49422 109200 49478 110000 6 o[58]
port 341 nsew signal output
rlabel metal2 s 50250 109200 50306 110000 6 o[59]
port 342 nsew signal output
rlabel metal2 s 4618 109200 4674 110000 6 o[5]
port 343 nsew signal output
rlabel metal2 s 51170 109200 51226 110000 6 o[60]
port 344 nsew signal output
rlabel metal2 s 51998 109200 52054 110000 6 o[61]
port 345 nsew signal output
rlabel metal2 s 52826 109200 52882 110000 6 o[62]
port 346 nsew signal output
rlabel metal2 s 53654 109200 53710 110000 6 o[63]
port 347 nsew signal output
rlabel metal2 s 54482 109200 54538 110000 6 o[64]
port 348 nsew signal output
rlabel metal2 s 55402 109200 55458 110000 6 o[65]
port 349 nsew signal output
rlabel metal2 s 56230 109200 56286 110000 6 o[66]
port 350 nsew signal output
rlabel metal2 s 57058 109200 57114 110000 6 o[67]
port 351 nsew signal output
rlabel metal2 s 57886 109200 57942 110000 6 o[68]
port 352 nsew signal output
rlabel metal2 s 58714 109200 58770 110000 6 o[69]
port 353 nsew signal output
rlabel metal2 s 5446 109200 5502 110000 6 o[6]
port 354 nsew signal output
rlabel metal2 s 59634 109200 59690 110000 6 o[70]
port 355 nsew signal output
rlabel metal2 s 60462 109200 60518 110000 6 o[71]
port 356 nsew signal output
rlabel metal2 s 61290 109200 61346 110000 6 o[72]
port 357 nsew signal output
rlabel metal2 s 62118 109200 62174 110000 6 o[73]
port 358 nsew signal output
rlabel metal2 s 62946 109200 63002 110000 6 o[74]
port 359 nsew signal output
rlabel metal2 s 63866 109200 63922 110000 6 o[75]
port 360 nsew signal output
rlabel metal2 s 64694 109200 64750 110000 6 o[76]
port 361 nsew signal output
rlabel metal2 s 65522 109200 65578 110000 6 o[77]
port 362 nsew signal output
rlabel metal2 s 66350 109200 66406 110000 6 o[78]
port 363 nsew signal output
rlabel metal2 s 67178 109200 67234 110000 6 o[79]
port 364 nsew signal output
rlabel metal2 s 6274 109200 6330 110000 6 o[7]
port 365 nsew signal output
rlabel metal2 s 68098 109200 68154 110000 6 o[80]
port 366 nsew signal output
rlabel metal2 s 68926 109200 68982 110000 6 o[81]
port 367 nsew signal output
rlabel metal2 s 69754 109200 69810 110000 6 o[82]
port 368 nsew signal output
rlabel metal2 s 70582 109200 70638 110000 6 o[83]
port 369 nsew signal output
rlabel metal2 s 71410 109200 71466 110000 6 o[84]
port 370 nsew signal output
rlabel metal2 s 72330 109200 72386 110000 6 o[85]
port 371 nsew signal output
rlabel metal2 s 73158 109200 73214 110000 6 o[86]
port 372 nsew signal output
rlabel metal2 s 73986 109200 74042 110000 6 o[87]
port 373 nsew signal output
rlabel metal2 s 74814 109200 74870 110000 6 o[88]
port 374 nsew signal output
rlabel metal2 s 75642 109200 75698 110000 6 o[89]
port 375 nsew signal output
rlabel metal2 s 7102 109200 7158 110000 6 o[8]
port 376 nsew signal output
rlabel metal2 s 76562 109200 76618 110000 6 o[90]
port 377 nsew signal output
rlabel metal2 s 77390 109200 77446 110000 6 o[91]
port 378 nsew signal output
rlabel metal2 s 78218 109200 78274 110000 6 o[92]
port 379 nsew signal output
rlabel metal2 s 79046 109200 79102 110000 6 o[93]
port 380 nsew signal output
rlabel metal2 s 79874 109200 79930 110000 6 o[94]
port 381 nsew signal output
rlabel metal2 s 80794 109200 80850 110000 6 o[95]
port 382 nsew signal output
rlabel metal2 s 81622 109200 81678 110000 6 o[96]
port 383 nsew signal output
rlabel metal2 s 82450 109200 82506 110000 6 o[97]
port 384 nsew signal output
rlabel metal2 s 83278 109200 83334 110000 6 o[98]
port 385 nsew signal output
rlabel metal2 s 84106 109200 84162 110000 6 o[99]
port 386 nsew signal output
rlabel metal2 s 7930 109200 7986 110000 6 o[9]
port 387 nsew signal output
rlabel metal2 s 108670 109200 108726 110000 6 rst
port 388 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32834300
string GDS_FILE /home/anton_unencrypted/shuttle-3/caravel_user_project/openlane/multiply_add_64x64/runs/multiply_add_64x64/results/finishing/multiply_add_64x64.magic.gds
string GDS_START 302210
<< end >>

