magic
tech sky130A
magscale 1 2
timestamp 1647885844
<< obsli1 >>
rect 1104 2159 228896 227409
<< obsm1 >>
rect 382 756 229894 227440
<< metal2 >>
rect 3790 229200 3846 230000
rect 11426 229200 11482 230000
rect 19062 229200 19118 230000
rect 26790 229200 26846 230000
rect 34426 229200 34482 230000
rect 42062 229200 42118 230000
rect 49790 229200 49846 230000
rect 57426 229200 57482 230000
rect 65062 229200 65118 230000
rect 72790 229200 72846 230000
rect 80426 229200 80482 230000
rect 88062 229200 88118 230000
rect 95790 229200 95846 230000
rect 103426 229200 103482 230000
rect 111062 229200 111118 230000
rect 118790 229200 118846 230000
rect 126426 229200 126482 230000
rect 134062 229200 134118 230000
rect 141790 229200 141846 230000
rect 149426 229200 149482 230000
rect 157062 229200 157118 230000
rect 164790 229200 164846 230000
rect 172426 229200 172482 230000
rect 180062 229200 180118 230000
rect 187790 229200 187846 230000
rect 195426 229200 195482 230000
rect 203062 229200 203118 230000
rect 210790 229200 210846 230000
rect 218426 229200 218482 230000
rect 226062 229200 226118 230000
rect 846 0 902 800
rect 2594 0 2650 800
rect 4434 0 4490 800
rect 6182 0 6238 800
rect 8022 0 8078 800
rect 9770 0 9826 800
rect 11610 0 11666 800
rect 13358 0 13414 800
rect 15198 0 15254 800
rect 16946 0 17002 800
rect 18786 0 18842 800
rect 20534 0 20590 800
rect 22374 0 22430 800
rect 24122 0 24178 800
rect 25962 0 26018 800
rect 27710 0 27766 800
rect 29550 0 29606 800
rect 31390 0 31446 800
rect 33138 0 33194 800
rect 34978 0 35034 800
rect 36726 0 36782 800
rect 38566 0 38622 800
rect 40314 0 40370 800
rect 42154 0 42210 800
rect 43902 0 43958 800
rect 45742 0 45798 800
rect 47490 0 47546 800
rect 49330 0 49386 800
rect 51078 0 51134 800
rect 52918 0 52974 800
rect 54666 0 54722 800
rect 56506 0 56562 800
rect 58346 0 58402 800
rect 60094 0 60150 800
rect 61934 0 61990 800
rect 63682 0 63738 800
rect 65522 0 65578 800
rect 67270 0 67326 800
rect 69110 0 69166 800
rect 70858 0 70914 800
rect 72698 0 72754 800
rect 74446 0 74502 800
rect 76286 0 76342 800
rect 78034 0 78090 800
rect 79874 0 79930 800
rect 81622 0 81678 800
rect 83462 0 83518 800
rect 85210 0 85266 800
rect 87050 0 87106 800
rect 88890 0 88946 800
rect 90638 0 90694 800
rect 92478 0 92534 800
rect 94226 0 94282 800
rect 96066 0 96122 800
rect 97814 0 97870 800
rect 99654 0 99710 800
rect 101402 0 101458 800
rect 103242 0 103298 800
rect 104990 0 105046 800
rect 106830 0 106886 800
rect 108578 0 108634 800
rect 110418 0 110474 800
rect 112166 0 112222 800
rect 114006 0 114062 800
rect 115846 0 115902 800
rect 117594 0 117650 800
rect 119434 0 119490 800
rect 121182 0 121238 800
rect 123022 0 123078 800
rect 124770 0 124826 800
rect 126610 0 126666 800
rect 128358 0 128414 800
rect 130198 0 130254 800
rect 131946 0 132002 800
rect 133786 0 133842 800
rect 135534 0 135590 800
rect 137374 0 137430 800
rect 139122 0 139178 800
rect 140962 0 141018 800
rect 142710 0 142766 800
rect 144550 0 144606 800
rect 146390 0 146446 800
rect 148138 0 148194 800
rect 149978 0 150034 800
rect 151726 0 151782 800
rect 153566 0 153622 800
rect 155314 0 155370 800
rect 157154 0 157210 800
rect 158902 0 158958 800
rect 160742 0 160798 800
rect 162490 0 162546 800
rect 164330 0 164386 800
rect 166078 0 166134 800
rect 167918 0 167974 800
rect 169666 0 169722 800
rect 171506 0 171562 800
rect 173346 0 173402 800
rect 175094 0 175150 800
rect 176934 0 176990 800
rect 178682 0 178738 800
rect 180522 0 180578 800
rect 182270 0 182326 800
rect 184110 0 184166 800
rect 185858 0 185914 800
rect 187698 0 187754 800
rect 189446 0 189502 800
rect 191286 0 191342 800
rect 193034 0 193090 800
rect 194874 0 194930 800
rect 196622 0 196678 800
rect 198462 0 198518 800
rect 200210 0 200266 800
rect 202050 0 202106 800
rect 203890 0 203946 800
rect 205638 0 205694 800
rect 207478 0 207534 800
rect 209226 0 209282 800
rect 211066 0 211122 800
rect 212814 0 212870 800
rect 214654 0 214710 800
rect 216402 0 216458 800
rect 218242 0 218298 800
rect 219990 0 220046 800
rect 221830 0 221886 800
rect 223578 0 223634 800
rect 225418 0 225474 800
rect 227166 0 227222 800
rect 229006 0 229062 800
<< obsm2 >>
rect 388 229144 3734 229242
rect 3902 229144 11370 229242
rect 11538 229144 19006 229242
rect 19174 229144 26734 229242
rect 26902 229144 34370 229242
rect 34538 229144 42006 229242
rect 42174 229144 49734 229242
rect 49902 229144 57370 229242
rect 57538 229144 65006 229242
rect 65174 229144 72734 229242
rect 72902 229144 80370 229242
rect 80538 229144 88006 229242
rect 88174 229144 95734 229242
rect 95902 229144 103370 229242
rect 103538 229144 111006 229242
rect 111174 229144 118734 229242
rect 118902 229144 126370 229242
rect 126538 229144 134006 229242
rect 134174 229144 141734 229242
rect 141902 229144 149370 229242
rect 149538 229144 157006 229242
rect 157174 229144 164734 229242
rect 164902 229144 172370 229242
rect 172538 229144 180006 229242
rect 180174 229144 187734 229242
rect 187902 229144 195370 229242
rect 195538 229144 203006 229242
rect 203174 229144 210734 229242
rect 210902 229144 218370 229242
rect 218538 229144 226006 229242
rect 226174 229144 229888 229242
rect 388 856 229888 229144
rect 388 734 790 856
rect 958 734 2538 856
rect 2706 734 4378 856
rect 4546 734 6126 856
rect 6294 734 7966 856
rect 8134 734 9714 856
rect 9882 734 11554 856
rect 11722 734 13302 856
rect 13470 734 15142 856
rect 15310 734 16890 856
rect 17058 734 18730 856
rect 18898 734 20478 856
rect 20646 734 22318 856
rect 22486 734 24066 856
rect 24234 734 25906 856
rect 26074 734 27654 856
rect 27822 734 29494 856
rect 29662 734 31334 856
rect 31502 734 33082 856
rect 33250 734 34922 856
rect 35090 734 36670 856
rect 36838 734 38510 856
rect 38678 734 40258 856
rect 40426 734 42098 856
rect 42266 734 43846 856
rect 44014 734 45686 856
rect 45854 734 47434 856
rect 47602 734 49274 856
rect 49442 734 51022 856
rect 51190 734 52862 856
rect 53030 734 54610 856
rect 54778 734 56450 856
rect 56618 734 58290 856
rect 58458 734 60038 856
rect 60206 734 61878 856
rect 62046 734 63626 856
rect 63794 734 65466 856
rect 65634 734 67214 856
rect 67382 734 69054 856
rect 69222 734 70802 856
rect 70970 734 72642 856
rect 72810 734 74390 856
rect 74558 734 76230 856
rect 76398 734 77978 856
rect 78146 734 79818 856
rect 79986 734 81566 856
rect 81734 734 83406 856
rect 83574 734 85154 856
rect 85322 734 86994 856
rect 87162 734 88834 856
rect 89002 734 90582 856
rect 90750 734 92422 856
rect 92590 734 94170 856
rect 94338 734 96010 856
rect 96178 734 97758 856
rect 97926 734 99598 856
rect 99766 734 101346 856
rect 101514 734 103186 856
rect 103354 734 104934 856
rect 105102 734 106774 856
rect 106942 734 108522 856
rect 108690 734 110362 856
rect 110530 734 112110 856
rect 112278 734 113950 856
rect 114118 734 115790 856
rect 115958 734 117538 856
rect 117706 734 119378 856
rect 119546 734 121126 856
rect 121294 734 122966 856
rect 123134 734 124714 856
rect 124882 734 126554 856
rect 126722 734 128302 856
rect 128470 734 130142 856
rect 130310 734 131890 856
rect 132058 734 133730 856
rect 133898 734 135478 856
rect 135646 734 137318 856
rect 137486 734 139066 856
rect 139234 734 140906 856
rect 141074 734 142654 856
rect 142822 734 144494 856
rect 144662 734 146334 856
rect 146502 734 148082 856
rect 148250 734 149922 856
rect 150090 734 151670 856
rect 151838 734 153510 856
rect 153678 734 155258 856
rect 155426 734 157098 856
rect 157266 734 158846 856
rect 159014 734 160686 856
rect 160854 734 162434 856
rect 162602 734 164274 856
rect 164442 734 166022 856
rect 166190 734 167862 856
rect 168030 734 169610 856
rect 169778 734 171450 856
rect 171618 734 173290 856
rect 173458 734 175038 856
rect 175206 734 176878 856
rect 177046 734 178626 856
rect 178794 734 180466 856
rect 180634 734 182214 856
rect 182382 734 184054 856
rect 184222 734 185802 856
rect 185970 734 187642 856
rect 187810 734 189390 856
rect 189558 734 191230 856
rect 191398 734 192978 856
rect 193146 734 194818 856
rect 194986 734 196566 856
rect 196734 734 198406 856
rect 198574 734 200154 856
rect 200322 734 201994 856
rect 202162 734 203834 856
rect 204002 734 205582 856
rect 205750 734 207422 856
rect 207590 734 209170 856
rect 209338 734 211010 856
rect 211178 734 212758 856
rect 212926 734 214598 856
rect 214766 734 216346 856
rect 216514 734 218186 856
rect 218354 734 219934 856
rect 220102 734 221774 856
rect 221942 734 223522 856
rect 223690 734 225362 856
rect 225530 734 227110 856
rect 227278 734 228950 856
rect 229118 734 229888 856
<< metal3 >>
rect 0 228896 800 229016
rect 0 227128 800 227248
rect 0 225360 800 225480
rect 0 223592 800 223712
rect 0 221688 800 221808
rect 0 219920 800 220040
rect 0 218152 800 218272
rect 0 216384 800 216504
rect 0 214616 800 214736
rect 0 212712 800 212832
rect 0 210944 800 211064
rect 0 209176 800 209296
rect 0 207408 800 207528
rect 0 205640 800 205760
rect 0 203736 800 203856
rect 0 201968 800 202088
rect 0 200200 800 200320
rect 0 198432 800 198552
rect 0 196528 800 196648
rect 0 194760 800 194880
rect 0 192992 800 193112
rect 0 191224 800 191344
rect 0 189456 800 189576
rect 0 187552 800 187672
rect 0 185784 800 185904
rect 0 184016 800 184136
rect 0 182248 800 182368
rect 0 180480 800 180600
rect 0 178576 800 178696
rect 0 176808 800 176928
rect 0 175040 800 175160
rect 0 173272 800 173392
rect 0 171504 800 171624
rect 0 169600 800 169720
rect 0 167832 800 167952
rect 0 166064 800 166184
rect 0 164296 800 164416
rect 0 162392 800 162512
rect 0 160624 800 160744
rect 0 158856 800 158976
rect 0 157088 800 157208
rect 0 155320 800 155440
rect 0 153416 800 153536
rect 0 151648 800 151768
rect 0 149880 800 150000
rect 0 148112 800 148232
rect 0 146344 800 146464
rect 0 144440 800 144560
rect 0 142672 800 142792
rect 0 140904 800 141024
rect 0 139136 800 139256
rect 0 137368 800 137488
rect 0 135464 800 135584
rect 0 133696 800 133816
rect 0 131928 800 132048
rect 0 130160 800 130280
rect 0 128256 800 128376
rect 0 126488 800 126608
rect 0 124720 800 124840
rect 0 122952 800 123072
rect 0 121184 800 121304
rect 0 119280 800 119400
rect 0 117512 800 117632
rect 0 115744 800 115864
rect 0 113976 800 114096
rect 0 112208 800 112328
rect 0 110304 800 110424
rect 0 108536 800 108656
rect 0 106768 800 106888
rect 0 105000 800 105120
rect 0 103232 800 103352
rect 0 101328 800 101448
rect 0 99560 800 99680
rect 0 97792 800 97912
rect 0 96024 800 96144
rect 0 94120 800 94240
rect 0 92352 800 92472
rect 0 90584 800 90704
rect 0 88816 800 88936
rect 0 87048 800 87168
rect 0 85144 800 85264
rect 0 83376 800 83496
rect 0 81608 800 81728
rect 0 79840 800 79960
rect 0 78072 800 78192
rect 0 76168 800 76288
rect 0 74400 800 74520
rect 0 72632 800 72752
rect 0 70864 800 70984
rect 0 69096 800 69216
rect 0 67192 800 67312
rect 0 65424 800 65544
rect 0 63656 800 63776
rect 0 61888 800 62008
rect 0 59984 800 60104
rect 0 58216 800 58336
rect 0 56448 800 56568
rect 0 54680 800 54800
rect 0 52912 800 53032
rect 0 51008 800 51128
rect 0 49240 800 49360
rect 0 47472 800 47592
rect 0 45704 800 45824
rect 0 43936 800 44056
rect 0 42032 800 42152
rect 0 40264 800 40384
rect 0 38496 800 38616
rect 0 36728 800 36848
rect 0 34960 800 35080
rect 0 33056 800 33176
rect 0 31288 800 31408
rect 0 29520 800 29640
rect 0 27752 800 27872
rect 0 25848 800 25968
rect 0 24080 800 24200
rect 0 22312 800 22432
rect 0 20544 800 20664
rect 0 18776 800 18896
rect 0 16872 800 16992
rect 0 15104 800 15224
rect 0 13336 800 13456
rect 0 11568 800 11688
rect 0 9800 800 9920
rect 0 7896 800 8016
rect 0 6128 800 6248
rect 0 4360 800 4480
rect 0 2592 800 2712
rect 0 824 800 944
<< obsm3 >>
rect 880 228816 229435 228989
rect 606 227328 229435 228816
rect 880 227048 229435 227328
rect 606 225560 229435 227048
rect 880 225280 229435 225560
rect 606 223792 229435 225280
rect 880 223512 229435 223792
rect 606 221888 229435 223512
rect 880 221608 229435 221888
rect 606 220120 229435 221608
rect 880 219840 229435 220120
rect 606 218352 229435 219840
rect 880 218072 229435 218352
rect 606 216584 229435 218072
rect 880 216304 229435 216584
rect 606 214816 229435 216304
rect 880 214536 229435 214816
rect 606 212912 229435 214536
rect 880 212632 229435 212912
rect 606 211144 229435 212632
rect 880 210864 229435 211144
rect 606 209376 229435 210864
rect 880 209096 229435 209376
rect 606 207608 229435 209096
rect 880 207328 229435 207608
rect 606 205840 229435 207328
rect 880 205560 229435 205840
rect 606 203936 229435 205560
rect 880 203656 229435 203936
rect 606 202168 229435 203656
rect 880 201888 229435 202168
rect 606 200400 229435 201888
rect 880 200120 229435 200400
rect 606 198632 229435 200120
rect 880 198352 229435 198632
rect 606 196728 229435 198352
rect 880 196448 229435 196728
rect 606 194960 229435 196448
rect 880 194680 229435 194960
rect 606 193192 229435 194680
rect 880 192912 229435 193192
rect 606 191424 229435 192912
rect 880 191144 229435 191424
rect 606 189656 229435 191144
rect 880 189376 229435 189656
rect 606 187752 229435 189376
rect 880 187472 229435 187752
rect 606 185984 229435 187472
rect 880 185704 229435 185984
rect 606 184216 229435 185704
rect 880 183936 229435 184216
rect 606 182448 229435 183936
rect 880 182168 229435 182448
rect 606 180680 229435 182168
rect 880 180400 229435 180680
rect 606 178776 229435 180400
rect 880 178496 229435 178776
rect 606 177008 229435 178496
rect 880 176728 229435 177008
rect 606 175240 229435 176728
rect 880 174960 229435 175240
rect 606 173472 229435 174960
rect 880 173192 229435 173472
rect 606 171704 229435 173192
rect 880 171424 229435 171704
rect 606 169800 229435 171424
rect 880 169520 229435 169800
rect 606 168032 229435 169520
rect 880 167752 229435 168032
rect 606 166264 229435 167752
rect 880 165984 229435 166264
rect 606 164496 229435 165984
rect 880 164216 229435 164496
rect 606 162592 229435 164216
rect 880 162312 229435 162592
rect 606 160824 229435 162312
rect 880 160544 229435 160824
rect 606 159056 229435 160544
rect 880 158776 229435 159056
rect 606 157288 229435 158776
rect 880 157008 229435 157288
rect 606 155520 229435 157008
rect 880 155240 229435 155520
rect 606 153616 229435 155240
rect 880 153336 229435 153616
rect 606 151848 229435 153336
rect 880 151568 229435 151848
rect 606 150080 229435 151568
rect 880 149800 229435 150080
rect 606 148312 229435 149800
rect 880 148032 229435 148312
rect 606 146544 229435 148032
rect 880 146264 229435 146544
rect 606 144640 229435 146264
rect 880 144360 229435 144640
rect 606 142872 229435 144360
rect 880 142592 229435 142872
rect 606 141104 229435 142592
rect 880 140824 229435 141104
rect 606 139336 229435 140824
rect 880 139056 229435 139336
rect 606 137568 229435 139056
rect 880 137288 229435 137568
rect 606 135664 229435 137288
rect 880 135384 229435 135664
rect 606 133896 229435 135384
rect 880 133616 229435 133896
rect 606 132128 229435 133616
rect 880 131848 229435 132128
rect 606 130360 229435 131848
rect 880 130080 229435 130360
rect 606 128456 229435 130080
rect 880 128176 229435 128456
rect 606 126688 229435 128176
rect 880 126408 229435 126688
rect 606 124920 229435 126408
rect 880 124640 229435 124920
rect 606 123152 229435 124640
rect 880 122872 229435 123152
rect 606 121384 229435 122872
rect 880 121104 229435 121384
rect 606 119480 229435 121104
rect 880 119200 229435 119480
rect 606 117712 229435 119200
rect 880 117432 229435 117712
rect 606 115944 229435 117432
rect 880 115664 229435 115944
rect 606 114176 229435 115664
rect 880 113896 229435 114176
rect 606 112408 229435 113896
rect 880 112128 229435 112408
rect 606 110504 229435 112128
rect 880 110224 229435 110504
rect 606 108736 229435 110224
rect 880 108456 229435 108736
rect 606 106968 229435 108456
rect 880 106688 229435 106968
rect 606 105200 229435 106688
rect 880 104920 229435 105200
rect 606 103432 229435 104920
rect 880 103152 229435 103432
rect 606 101528 229435 103152
rect 880 101248 229435 101528
rect 606 99760 229435 101248
rect 880 99480 229435 99760
rect 606 97992 229435 99480
rect 880 97712 229435 97992
rect 606 96224 229435 97712
rect 880 95944 229435 96224
rect 606 94320 229435 95944
rect 880 94040 229435 94320
rect 606 92552 229435 94040
rect 880 92272 229435 92552
rect 606 90784 229435 92272
rect 880 90504 229435 90784
rect 606 89016 229435 90504
rect 880 88736 229435 89016
rect 606 87248 229435 88736
rect 880 86968 229435 87248
rect 606 85344 229435 86968
rect 880 85064 229435 85344
rect 606 83576 229435 85064
rect 880 83296 229435 83576
rect 606 81808 229435 83296
rect 880 81528 229435 81808
rect 606 80040 229435 81528
rect 880 79760 229435 80040
rect 606 78272 229435 79760
rect 880 77992 229435 78272
rect 606 76368 229435 77992
rect 880 76088 229435 76368
rect 606 74600 229435 76088
rect 880 74320 229435 74600
rect 606 72832 229435 74320
rect 880 72552 229435 72832
rect 606 71064 229435 72552
rect 880 70784 229435 71064
rect 606 69296 229435 70784
rect 880 69016 229435 69296
rect 606 67392 229435 69016
rect 880 67112 229435 67392
rect 606 65624 229435 67112
rect 880 65344 229435 65624
rect 606 63856 229435 65344
rect 880 63576 229435 63856
rect 606 62088 229435 63576
rect 880 61808 229435 62088
rect 606 60184 229435 61808
rect 880 59904 229435 60184
rect 606 58416 229435 59904
rect 880 58136 229435 58416
rect 606 56648 229435 58136
rect 880 56368 229435 56648
rect 606 54880 229435 56368
rect 880 54600 229435 54880
rect 606 53112 229435 54600
rect 880 52832 229435 53112
rect 606 51208 229435 52832
rect 880 50928 229435 51208
rect 606 49440 229435 50928
rect 880 49160 229435 49440
rect 606 47672 229435 49160
rect 880 47392 229435 47672
rect 606 45904 229435 47392
rect 880 45624 229435 45904
rect 606 44136 229435 45624
rect 880 43856 229435 44136
rect 606 42232 229435 43856
rect 880 41952 229435 42232
rect 606 40464 229435 41952
rect 880 40184 229435 40464
rect 606 38696 229435 40184
rect 880 38416 229435 38696
rect 606 36928 229435 38416
rect 880 36648 229435 36928
rect 606 35160 229435 36648
rect 880 34880 229435 35160
rect 606 33256 229435 34880
rect 880 32976 229435 33256
rect 606 31488 229435 32976
rect 880 31208 229435 31488
rect 606 29720 229435 31208
rect 880 29440 229435 29720
rect 606 27952 229435 29440
rect 880 27672 229435 27952
rect 606 26048 229435 27672
rect 880 25768 229435 26048
rect 606 24280 229435 25768
rect 880 24000 229435 24280
rect 606 22512 229435 24000
rect 880 22232 229435 22512
rect 606 20744 229435 22232
rect 880 20464 229435 20744
rect 606 18976 229435 20464
rect 880 18696 229435 18976
rect 606 17072 229435 18696
rect 880 16792 229435 17072
rect 606 15304 229435 16792
rect 880 15024 229435 15304
rect 606 13536 229435 15024
rect 880 13256 229435 13536
rect 606 11768 229435 13256
rect 880 11488 229435 11768
rect 606 10000 229435 11488
rect 880 9720 229435 10000
rect 606 8096 229435 9720
rect 880 7816 229435 8096
rect 606 6328 229435 7816
rect 880 6048 229435 6328
rect 606 4560 229435 6048
rect 880 4280 229435 4560
rect 606 2792 229435 4280
rect 880 2512 229435 2792
rect 606 1024 229435 2512
rect 880 851 229435 1024
<< metal4 >>
rect 1794 2128 2414 227440
rect 19794 2128 20414 227440
rect 37794 2128 38414 227440
rect 55794 2128 56414 227440
rect 73794 2128 74414 227440
rect 91794 2128 92414 227440
rect 109794 2128 110414 227440
rect 127794 2128 128414 227440
rect 145794 2128 146414 227440
rect 163794 2128 164414 227440
rect 181794 2128 182414 227440
rect 199794 2128 200414 227440
rect 217794 2128 218414 227440
<< obsm4 >>
rect 611 227520 227181 227629
rect 611 2048 1714 227520
rect 2494 2048 19714 227520
rect 20494 2048 37714 227520
rect 38494 2048 55714 227520
rect 56494 2048 73714 227520
rect 74494 2048 91714 227520
rect 92494 2048 109714 227520
rect 110494 2048 127714 227520
rect 128494 2048 145714 227520
rect 146494 2048 163714 227520
rect 164494 2048 181714 227520
rect 182494 2048 199714 227520
rect 200494 2048 217714 227520
rect 218494 2048 227181 227520
rect 611 1667 227181 2048
<< labels >>
rlabel metal2 s 3790 229200 3846 230000 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 824 800 944 6 D1[0]
port 2 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 D1[10]
port 3 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 D1[11]
port 4 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 D1[12]
port 5 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 D1[13]
port 6 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 D1[14]
port 7 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 D1[15]
port 8 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 D1[16]
port 9 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 D1[17]
port 10 nsew signal output
rlabel metal3 s 0 33056 800 33176 6 D1[18]
port 11 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 D1[19]
port 12 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 D1[1]
port 13 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 D1[20]
port 14 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 D1[21]
port 15 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 D1[22]
port 16 nsew signal output
rlabel metal3 s 0 42032 800 42152 6 D1[23]
port 17 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 D1[24]
port 18 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 D1[25]
port 19 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 D1[26]
port 20 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 D1[27]
port 21 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 D1[28]
port 22 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 D1[29]
port 23 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 D1[2]
port 24 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 D1[30]
port 25 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 D1[31]
port 26 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 D1[32]
port 27 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 D1[33]
port 28 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 D1[34]
port 29 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 D1[35]
port 30 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 D1[36]
port 31 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 D1[37]
port 32 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 D1[38]
port 33 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 D1[39]
port 34 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 D1[3]
port 35 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 D1[40]
port 36 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 D1[41]
port 37 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 D1[42]
port 38 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 D1[43]
port 39 nsew signal output
rlabel metal3 s 0 79840 800 79960 6 D1[44]
port 40 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 D1[45]
port 41 nsew signal output
rlabel metal3 s 0 83376 800 83496 6 D1[46]
port 42 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 D1[47]
port 43 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 D1[48]
port 44 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 D1[49]
port 45 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 D1[4]
port 46 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 D1[50]
port 47 nsew signal output
rlabel metal3 s 0 92352 800 92472 6 D1[51]
port 48 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 D1[52]
port 49 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 D1[53]
port 50 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 D1[54]
port 51 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 D1[55]
port 52 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 D1[56]
port 53 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 D1[57]
port 54 nsew signal output
rlabel metal3 s 0 105000 800 105120 6 D1[58]
port 55 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 D1[59]
port 56 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 D1[5]
port 57 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 D1[60]
port 58 nsew signal output
rlabel metal3 s 0 110304 800 110424 6 D1[61]
port 59 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 D1[62]
port 60 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 D1[63]
port 61 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 D1[6]
port 62 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 D1[7]
port 63 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 D1[8]
port 64 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 D1[9]
port 65 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 D2[0]
port 66 nsew signal output
rlabel metal3 s 0 133696 800 133816 6 D2[10]
port 67 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 D2[11]
port 68 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 D2[12]
port 69 nsew signal output
rlabel metal3 s 0 139136 800 139256 6 D2[13]
port 70 nsew signal output
rlabel metal3 s 0 140904 800 141024 6 D2[14]
port 71 nsew signal output
rlabel metal3 s 0 142672 800 142792 6 D2[15]
port 72 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 D2[16]
port 73 nsew signal output
rlabel metal3 s 0 146344 800 146464 6 D2[17]
port 74 nsew signal output
rlabel metal3 s 0 148112 800 148232 6 D2[18]
port 75 nsew signal output
rlabel metal3 s 0 149880 800 150000 6 D2[19]
port 76 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 D2[1]
port 77 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 D2[20]
port 78 nsew signal output
rlabel metal3 s 0 153416 800 153536 6 D2[21]
port 79 nsew signal output
rlabel metal3 s 0 155320 800 155440 6 D2[22]
port 80 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 D2[23]
port 81 nsew signal output
rlabel metal3 s 0 158856 800 158976 6 D2[24]
port 82 nsew signal output
rlabel metal3 s 0 160624 800 160744 6 D2[25]
port 83 nsew signal output
rlabel metal3 s 0 162392 800 162512 6 D2[26]
port 84 nsew signal output
rlabel metal3 s 0 164296 800 164416 6 D2[27]
port 85 nsew signal output
rlabel metal3 s 0 166064 800 166184 6 D2[28]
port 86 nsew signal output
rlabel metal3 s 0 167832 800 167952 6 D2[29]
port 87 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 D2[2]
port 88 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 D2[30]
port 89 nsew signal output
rlabel metal3 s 0 171504 800 171624 6 D2[31]
port 90 nsew signal output
rlabel metal3 s 0 173272 800 173392 6 D2[32]
port 91 nsew signal output
rlabel metal3 s 0 175040 800 175160 6 D2[33]
port 92 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 D2[34]
port 93 nsew signal output
rlabel metal3 s 0 178576 800 178696 6 D2[35]
port 94 nsew signal output
rlabel metal3 s 0 180480 800 180600 6 D2[36]
port 95 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 D2[37]
port 96 nsew signal output
rlabel metal3 s 0 184016 800 184136 6 D2[38]
port 97 nsew signal output
rlabel metal3 s 0 185784 800 185904 6 D2[39]
port 98 nsew signal output
rlabel metal3 s 0 121184 800 121304 6 D2[3]
port 99 nsew signal output
rlabel metal3 s 0 187552 800 187672 6 D2[40]
port 100 nsew signal output
rlabel metal3 s 0 189456 800 189576 6 D2[41]
port 101 nsew signal output
rlabel metal3 s 0 191224 800 191344 6 D2[42]
port 102 nsew signal output
rlabel metal3 s 0 192992 800 193112 6 D2[43]
port 103 nsew signal output
rlabel metal3 s 0 194760 800 194880 6 D2[44]
port 104 nsew signal output
rlabel metal3 s 0 196528 800 196648 6 D2[45]
port 105 nsew signal output
rlabel metal3 s 0 198432 800 198552 6 D2[46]
port 106 nsew signal output
rlabel metal3 s 0 200200 800 200320 6 D2[47]
port 107 nsew signal output
rlabel metal3 s 0 201968 800 202088 6 D2[48]
port 108 nsew signal output
rlabel metal3 s 0 203736 800 203856 6 D2[49]
port 109 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 D2[4]
port 110 nsew signal output
rlabel metal3 s 0 205640 800 205760 6 D2[50]
port 111 nsew signal output
rlabel metal3 s 0 207408 800 207528 6 D2[51]
port 112 nsew signal output
rlabel metal3 s 0 209176 800 209296 6 D2[52]
port 113 nsew signal output
rlabel metal3 s 0 210944 800 211064 6 D2[53]
port 114 nsew signal output
rlabel metal3 s 0 212712 800 212832 6 D2[54]
port 115 nsew signal output
rlabel metal3 s 0 214616 800 214736 6 D2[55]
port 116 nsew signal output
rlabel metal3 s 0 216384 800 216504 6 D2[56]
port 117 nsew signal output
rlabel metal3 s 0 218152 800 218272 6 D2[57]
port 118 nsew signal output
rlabel metal3 s 0 219920 800 220040 6 D2[58]
port 119 nsew signal output
rlabel metal3 s 0 221688 800 221808 6 D2[59]
port 120 nsew signal output
rlabel metal3 s 0 124720 800 124840 6 D2[5]
port 121 nsew signal output
rlabel metal3 s 0 223592 800 223712 6 D2[60]
port 122 nsew signal output
rlabel metal3 s 0 225360 800 225480 6 D2[61]
port 123 nsew signal output
rlabel metal3 s 0 227128 800 227248 6 D2[62]
port 124 nsew signal output
rlabel metal3 s 0 228896 800 229016 6 D2[63]
port 125 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 D2[6]
port 126 nsew signal output
rlabel metal3 s 0 128256 800 128376 6 D2[7]
port 127 nsew signal output
rlabel metal3 s 0 130160 800 130280 6 D2[8]
port 128 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 D2[9]
port 129 nsew signal output
rlabel metal2 s 846 0 902 800 6 D3[0]
port 130 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 D3[10]
port 131 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 D3[11]
port 132 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 D3[12]
port 133 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 D3[13]
port 134 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 D3[14]
port 135 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 D3[15]
port 136 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 D3[16]
port 137 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 D3[17]
port 138 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 D3[18]
port 139 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 D3[19]
port 140 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 D3[1]
port 141 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 D3[20]
port 142 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 D3[21]
port 143 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 D3[22]
port 144 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 D3[23]
port 145 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 D3[24]
port 146 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 D3[25]
port 147 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 D3[26]
port 148 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 D3[27]
port 149 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 D3[28]
port 150 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 D3[29]
port 151 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 D3[2]
port 152 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 D3[30]
port 153 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 D3[31]
port 154 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 D3[32]
port 155 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 D3[33]
port 156 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 D3[34]
port 157 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 D3[35]
port 158 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 D3[36]
port 159 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 D3[37]
port 160 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 D3[38]
port 161 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 D3[39]
port 162 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 D3[3]
port 163 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 D3[40]
port 164 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 D3[41]
port 165 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 D3[42]
port 166 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 D3[43]
port 167 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 D3[44]
port 168 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 D3[45]
port 169 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 D3[46]
port 170 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 D3[47]
port 171 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 D3[48]
port 172 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 D3[49]
port 173 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 D3[4]
port 174 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 D3[50]
port 175 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 D3[51]
port 176 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 D3[52]
port 177 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 D3[53]
port 178 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 D3[54]
port 179 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 D3[55]
port 180 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 D3[56]
port 181 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 D3[57]
port 182 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 D3[58]
port 183 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 D3[59]
port 184 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 D3[5]
port 185 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 D3[60]
port 186 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 D3[61]
port 187 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 D3[62]
port 188 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 D3[63]
port 189 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 D3[6]
port 190 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 D3[7]
port 191 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 D3[8]
port 192 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 D3[9]
port 193 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 DW[0]
port 194 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 DW[10]
port 195 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 DW[11]
port 196 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 DW[12]
port 197 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 DW[13]
port 198 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 DW[14]
port 199 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 DW[15]
port 200 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 DW[16]
port 201 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 DW[17]
port 202 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 DW[18]
port 203 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 DW[19]
port 204 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 DW[1]
port 205 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 DW[20]
port 206 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 DW[21]
port 207 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 DW[22]
port 208 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 DW[23]
port 209 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 DW[24]
port 210 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 DW[25]
port 211 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 DW[26]
port 212 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 DW[27]
port 213 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 DW[28]
port 214 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 DW[29]
port 215 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 DW[2]
port 216 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 DW[30]
port 217 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 DW[31]
port 218 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 DW[32]
port 219 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 DW[33]
port 220 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 DW[34]
port 221 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 DW[35]
port 222 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 DW[36]
port 223 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 DW[37]
port 224 nsew signal input
rlabel metal2 s 184110 0 184166 800 6 DW[38]
port 225 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 DW[39]
port 226 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 DW[3]
port 227 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 DW[40]
port 228 nsew signal input
rlabel metal2 s 189446 0 189502 800 6 DW[41]
port 229 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 DW[42]
port 230 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 DW[43]
port 231 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 DW[44]
port 232 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 DW[45]
port 233 nsew signal input
rlabel metal2 s 198462 0 198518 800 6 DW[46]
port 234 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 DW[47]
port 235 nsew signal input
rlabel metal2 s 202050 0 202106 800 6 DW[48]
port 236 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 DW[49]
port 237 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 DW[4]
port 238 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 DW[50]
port 239 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 DW[51]
port 240 nsew signal input
rlabel metal2 s 209226 0 209282 800 6 DW[52]
port 241 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 DW[53]
port 242 nsew signal input
rlabel metal2 s 212814 0 212870 800 6 DW[54]
port 243 nsew signal input
rlabel metal2 s 214654 0 214710 800 6 DW[55]
port 244 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 DW[56]
port 245 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 DW[57]
port 246 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 DW[58]
port 247 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 DW[59]
port 248 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 DW[5]
port 249 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 DW[60]
port 250 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 DW[61]
port 251 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 DW[62]
port 252 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 DW[63]
port 253 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 DW[6]
port 254 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 DW[7]
port 255 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 DW[8]
port 256 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 DW[9]
port 257 nsew signal input
rlabel metal2 s 19062 229200 19118 230000 6 R1[0]
port 258 nsew signal input
rlabel metal2 s 26790 229200 26846 230000 6 R1[1]
port 259 nsew signal input
rlabel metal2 s 34426 229200 34482 230000 6 R1[2]
port 260 nsew signal input
rlabel metal2 s 42062 229200 42118 230000 6 R1[3]
port 261 nsew signal input
rlabel metal2 s 49790 229200 49846 230000 6 R1[4]
port 262 nsew signal input
rlabel metal2 s 57426 229200 57482 230000 6 R1[5]
port 263 nsew signal input
rlabel metal2 s 65062 229200 65118 230000 6 R1[6]
port 264 nsew signal input
rlabel metal2 s 72790 229200 72846 230000 6 R2[0]
port 265 nsew signal input
rlabel metal2 s 80426 229200 80482 230000 6 R2[1]
port 266 nsew signal input
rlabel metal2 s 88062 229200 88118 230000 6 R2[2]
port 267 nsew signal input
rlabel metal2 s 95790 229200 95846 230000 6 R2[3]
port 268 nsew signal input
rlabel metal2 s 103426 229200 103482 230000 6 R2[4]
port 269 nsew signal input
rlabel metal2 s 111062 229200 111118 230000 6 R2[5]
port 270 nsew signal input
rlabel metal2 s 118790 229200 118846 230000 6 R2[6]
port 271 nsew signal input
rlabel metal2 s 126426 229200 126482 230000 6 R3[0]
port 272 nsew signal input
rlabel metal2 s 134062 229200 134118 230000 6 R3[1]
port 273 nsew signal input
rlabel metal2 s 141790 229200 141846 230000 6 R3[2]
port 274 nsew signal input
rlabel metal2 s 149426 229200 149482 230000 6 R3[3]
port 275 nsew signal input
rlabel metal2 s 157062 229200 157118 230000 6 R3[4]
port 276 nsew signal input
rlabel metal2 s 164790 229200 164846 230000 6 R3[5]
port 277 nsew signal input
rlabel metal2 s 172426 229200 172482 230000 6 R3[6]
port 278 nsew signal input
rlabel metal2 s 180062 229200 180118 230000 6 RW[0]
port 279 nsew signal input
rlabel metal2 s 187790 229200 187846 230000 6 RW[1]
port 280 nsew signal input
rlabel metal2 s 195426 229200 195482 230000 6 RW[2]
port 281 nsew signal input
rlabel metal2 s 203062 229200 203118 230000 6 RW[3]
port 282 nsew signal input
rlabel metal2 s 210790 229200 210846 230000 6 RW[4]
port 283 nsew signal input
rlabel metal2 s 218426 229200 218482 230000 6 RW[5]
port 284 nsew signal input
rlabel metal2 s 226062 229200 226118 230000 6 RW[6]
port 285 nsew signal input
rlabel metal4 s 19794 2128 20414 227440 6 VGND
port 286 nsew ground input
rlabel metal4 s 55794 2128 56414 227440 6 VGND
port 286 nsew ground input
rlabel metal4 s 91794 2128 92414 227440 6 VGND
port 286 nsew ground input
rlabel metal4 s 127794 2128 128414 227440 6 VGND
port 286 nsew ground input
rlabel metal4 s 163794 2128 164414 227440 6 VGND
port 286 nsew ground input
rlabel metal4 s 199794 2128 200414 227440 6 VGND
port 286 nsew ground input
rlabel metal4 s 1794 2128 2414 227440 6 VPWR
port 287 nsew power input
rlabel metal4 s 37794 2128 38414 227440 6 VPWR
port 287 nsew power input
rlabel metal4 s 73794 2128 74414 227440 6 VPWR
port 287 nsew power input
rlabel metal4 s 109794 2128 110414 227440 6 VPWR
port 287 nsew power input
rlabel metal4 s 145794 2128 146414 227440 6 VPWR
port 287 nsew power input
rlabel metal4 s 181794 2128 182414 227440 6 VPWR
port 287 nsew power input
rlabel metal4 s 217794 2128 218414 227440 6 VPWR
port 287 nsew power input
rlabel metal2 s 11426 229200 11482 230000 6 WE
port 288 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 230000 230000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 115795734
string GDS_FILE /home/anton_unencrypted/shuttle-3/caravel_user_project/openlane/Microwatt_FP_DFFRFile/runs/Microwatt_FP_DFFRFile/results/finishing/Microwatt_FP_DFFRFile.magic.gds
string GDS_START 624536
<< end >>

