VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Microwatt_FP_DFFRFile
  CLASS BLOCK ;
  FOREIGN Microwatt_FP_DFFRFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 1150.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 1146.000 19.230 1150.000 ;
    END
  END CLK
  PIN D1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END D1[31]
  PIN D1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END D1[32]
  PIN D1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END D1[33]
  PIN D1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END D1[34]
  PIN D1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END D1[35]
  PIN D1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END D1[36]
  PIN D1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END D1[37]
  PIN D1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END D1[38]
  PIN D1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END D1[39]
  PIN D1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END D1[3]
  PIN D1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END D1[40]
  PIN D1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END D1[41]
  PIN D1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END D1[42]
  PIN D1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END D1[43]
  PIN D1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END D1[44]
  PIN D1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END D1[45]
  PIN D1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END D1[46]
  PIN D1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END D1[47]
  PIN D1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END D1[48]
  PIN D1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END D1[49]
  PIN D1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END D1[4]
  PIN D1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END D1[50]
  PIN D1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END D1[51]
  PIN D1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END D1[52]
  PIN D1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END D1[53]
  PIN D1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END D1[54]
  PIN D1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END D1[55]
  PIN D1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END D1[56]
  PIN D1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END D1[57]
  PIN D1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END D1[58]
  PIN D1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END D1[59]
  PIN D1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END D1[5]
  PIN D1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END D1[60]
  PIN D1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END D1[61]
  PIN D1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END D1[62]
  PIN D1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END D1[63]
  PIN D1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 4.000 741.160 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 830.320 4.000 830.920 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 857.520 4.000 858.120 ;
    END
  END D2[31]
  PIN D2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END D2[32]
  PIN D2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 4.000 875.800 ;
    END
  END D2[33]
  PIN D2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END D2[34]
  PIN D2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END D2[35]
  PIN D2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END D2[36]
  PIN D2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END D2[37]
  PIN D2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END D2[38]
  PIN D2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.920 4.000 929.520 ;
    END
  END D2[39]
  PIN D2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END D2[3]
  PIN D2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END D2[40]
  PIN D2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END D2[41]
  PIN D2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.120 4.000 956.720 ;
    END
  END D2[42]
  PIN D2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.960 4.000 965.560 ;
    END
  END D2[43]
  PIN D2[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.800 4.000 974.400 ;
    END
  END D2[44]
  PIN D2[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END D2[45]
  PIN D2[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END D2[46]
  PIN D2[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.000 4.000 1001.600 ;
    END
  END D2[47]
  PIN D2[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END D2[48]
  PIN D2[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END D2[49]
  PIN D2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END D2[4]
  PIN D2[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1028.200 4.000 1028.800 ;
    END
  END D2[50]
  PIN D2[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END D2[51]
  PIN D2[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.880 4.000 1046.480 ;
    END
  END D2[52]
  PIN D2[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.720 4.000 1055.320 ;
    END
  END D2[53]
  PIN D2[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1063.560 4.000 1064.160 ;
    END
  END D2[54]
  PIN D2[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.080 4.000 1073.680 ;
    END
  END D2[55]
  PIN D2[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.920 4.000 1082.520 ;
    END
  END D2[56]
  PIN D2[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.760 4.000 1091.360 ;
    END
  END D2[57]
  PIN D2[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END D2[58]
  PIN D2[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END D2[59]
  PIN D2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END D2[5]
  PIN D2[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.960 4.000 1118.560 ;
    END
  END D2[60]
  PIN D2[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1126.800 4.000 1127.400 ;
    END
  END D2[61]
  PIN D2[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END D2[62]
  PIN D2[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1144.480 4.000 1145.080 ;
    END
  END D2[63]
  PIN D2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END D2[9]
  PIN D3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END D3[0]
  PIN D3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END D3[10]
  PIN D3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END D3[11]
  PIN D3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END D3[12]
  PIN D3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END D3[13]
  PIN D3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END D3[14]
  PIN D3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END D3[15]
  PIN D3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END D3[16]
  PIN D3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END D3[17]
  PIN D3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END D3[18]
  PIN D3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END D3[19]
  PIN D3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END D3[1]
  PIN D3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END D3[20]
  PIN D3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END D3[21]
  PIN D3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END D3[22]
  PIN D3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END D3[23]
  PIN D3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END D3[24]
  PIN D3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END D3[25]
  PIN D3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END D3[26]
  PIN D3[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END D3[27]
  PIN D3[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END D3[28]
  PIN D3[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END D3[29]
  PIN D3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END D3[2]
  PIN D3[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END D3[30]
  PIN D3[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END D3[31]
  PIN D3[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END D3[32]
  PIN D3[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END D3[33]
  PIN D3[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END D3[34]
  PIN D3[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END D3[35]
  PIN D3[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END D3[36]
  PIN D3[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END D3[37]
  PIN D3[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END D3[38]
  PIN D3[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END D3[39]
  PIN D3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END D3[3]
  PIN D3[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END D3[40]
  PIN D3[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END D3[41]
  PIN D3[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END D3[42]
  PIN D3[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END D3[43]
  PIN D3[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END D3[44]
  PIN D3[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END D3[45]
  PIN D3[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END D3[46]
  PIN D3[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END D3[47]
  PIN D3[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END D3[48]
  PIN D3[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END D3[49]
  PIN D3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END D3[4]
  PIN D3[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END D3[50]
  PIN D3[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END D3[51]
  PIN D3[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END D3[52]
  PIN D3[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END D3[53]
  PIN D3[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END D3[54]
  PIN D3[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END D3[55]
  PIN D3[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END D3[56]
  PIN D3[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END D3[57]
  PIN D3[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END D3[58]
  PIN D3[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END D3[59]
  PIN D3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END D3[5]
  PIN D3[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END D3[60]
  PIN D3[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END D3[61]
  PIN D3[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END D3[62]
  PIN D3[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END D3[63]
  PIN D3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END D3[6]
  PIN D3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END D3[7]
  PIN D3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END D3[8]
  PIN D3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END D3[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 0.000 768.110 4.000 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 0.000 803.990 4.000 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 0.000 857.810 4.000 ;
    END
  END DW[31]
  PIN DW[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END DW[32]
  PIN DW[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 0.000 875.750 4.000 ;
    END
  END DW[33]
  PIN DW[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 4.000 ;
    END
  END DW[34]
  PIN DW[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END DW[35]
  PIN DW[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END DW[36]
  PIN DW[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END DW[37]
  PIN DW[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END DW[38]
  PIN DW[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END DW[39]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END DW[3]
  PIN DW[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END DW[40]
  PIN DW[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END DW[41]
  PIN DW[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END DW[42]
  PIN DW[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END DW[43]
  PIN DW[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 0.000 974.650 4.000 ;
    END
  END DW[44]
  PIN DW[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END DW[45]
  PIN DW[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END DW[46]
  PIN DW[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.050 0.000 1001.330 4.000 ;
    END
  END DW[47]
  PIN DW[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 0.000 1010.530 4.000 ;
    END
  END DW[48]
  PIN DW[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.450 0.000 1019.730 4.000 ;
    END
  END DW[49]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END DW[4]
  PIN DW[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.190 0.000 1028.470 4.000 ;
    END
  END DW[50]
  PIN DW[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END DW[51]
  PIN DW[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END DW[52]
  PIN DW[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END DW[53]
  PIN DW[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 0.000 1064.350 4.000 ;
    END
  END DW[54]
  PIN DW[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END DW[55]
  PIN DW[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END DW[56]
  PIN DW[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END DW[57]
  PIN DW[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 0.000 1100.230 4.000 ;
    END
  END DW[58]
  PIN DW[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END DW[59]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END DW[5]
  PIN DW[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 0.000 1118.170 4.000 ;
    END
  END DW[60]
  PIN DW[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END DW[61]
  PIN DW[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.830 0.000 1136.110 4.000 ;
    END
  END DW[62]
  PIN DW[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END DW[63]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END DW[9]
  PIN R1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 1146.000 95.590 1150.000 ;
    END
  END R1[0]
  PIN R1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 1146.000 134.230 1150.000 ;
    END
  END R1[1]
  PIN R1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 1146.000 172.410 1150.000 ;
    END
  END R1[2]
  PIN R1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 1146.000 210.590 1150.000 ;
    END
  END R1[3]
  PIN R1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 1146.000 249.230 1150.000 ;
    END
  END R1[4]
  PIN R1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 1146.000 287.410 1150.000 ;
    END
  END R1[5]
  PIN R1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1146.000 325.590 1150.000 ;
    END
  END R1[6]
  PIN R2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1146.000 364.230 1150.000 ;
    END
  END R2[0]
  PIN R2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 1146.000 402.410 1150.000 ;
    END
  END R2[1]
  PIN R2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 1146.000 440.590 1150.000 ;
    END
  END R2[2]
  PIN R2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 1146.000 479.230 1150.000 ;
    END
  END R2[3]
  PIN R2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 1146.000 517.410 1150.000 ;
    END
  END R2[4]
  PIN R2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 1146.000 555.590 1150.000 ;
    END
  END R2[5]
  PIN R2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1146.000 594.230 1150.000 ;
    END
  END R2[6]
  PIN R3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 1146.000 632.410 1150.000 ;
    END
  END R3[0]
  PIN R3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 1146.000 670.590 1150.000 ;
    END
  END R3[1]
  PIN R3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 1146.000 709.230 1150.000 ;
    END
  END R3[2]
  PIN R3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1146.000 747.410 1150.000 ;
    END
  END R3[3]
  PIN R3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 1146.000 785.590 1150.000 ;
    END
  END R3[4]
  PIN R3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 1146.000 824.230 1150.000 ;
    END
  END R3[5]
  PIN R3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 1146.000 862.410 1150.000 ;
    END
  END R3[6]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 1146.000 900.590 1150.000 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 1146.000 939.230 1150.000 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 1146.000 977.410 1150.000 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 1146.000 1015.590 1150.000 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 1146.000 1054.230 1150.000 ;
    END
  END RW[4]
  PIN RW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 1146.000 1092.410 1150.000 ;
    END
  END RW[5]
  PIN RW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 1146.000 1130.590 1150.000 ;
    END
  END RW[6]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 10.640 642.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 10.640 822.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 10.640 1002.070 1137.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 10.640 912.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 1137.200 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 1146.000 57.410 1150.000 ;
    END
  END WE
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1144.480 1137.045 ;
      LAYER met1 ;
        RECT 1.910 3.780 1149.470 1137.200 ;
      LAYER met2 ;
        RECT 1.940 1145.720 18.670 1146.210 ;
        RECT 19.510 1145.720 56.850 1146.210 ;
        RECT 57.690 1145.720 95.030 1146.210 ;
        RECT 95.870 1145.720 133.670 1146.210 ;
        RECT 134.510 1145.720 171.850 1146.210 ;
        RECT 172.690 1145.720 210.030 1146.210 ;
        RECT 210.870 1145.720 248.670 1146.210 ;
        RECT 249.510 1145.720 286.850 1146.210 ;
        RECT 287.690 1145.720 325.030 1146.210 ;
        RECT 325.870 1145.720 363.670 1146.210 ;
        RECT 364.510 1145.720 401.850 1146.210 ;
        RECT 402.690 1145.720 440.030 1146.210 ;
        RECT 440.870 1145.720 478.670 1146.210 ;
        RECT 479.510 1145.720 516.850 1146.210 ;
        RECT 517.690 1145.720 555.030 1146.210 ;
        RECT 555.870 1145.720 593.670 1146.210 ;
        RECT 594.510 1145.720 631.850 1146.210 ;
        RECT 632.690 1145.720 670.030 1146.210 ;
        RECT 670.870 1145.720 708.670 1146.210 ;
        RECT 709.510 1145.720 746.850 1146.210 ;
        RECT 747.690 1145.720 785.030 1146.210 ;
        RECT 785.870 1145.720 823.670 1146.210 ;
        RECT 824.510 1145.720 861.850 1146.210 ;
        RECT 862.690 1145.720 900.030 1146.210 ;
        RECT 900.870 1145.720 938.670 1146.210 ;
        RECT 939.510 1145.720 976.850 1146.210 ;
        RECT 977.690 1145.720 1015.030 1146.210 ;
        RECT 1015.870 1145.720 1053.670 1146.210 ;
        RECT 1054.510 1145.720 1091.850 1146.210 ;
        RECT 1092.690 1145.720 1130.030 1146.210 ;
        RECT 1130.870 1145.720 1149.440 1146.210 ;
        RECT 1.940 4.280 1149.440 1145.720 ;
        RECT 1.940 3.670 3.950 4.280 ;
        RECT 4.790 3.670 12.690 4.280 ;
        RECT 13.530 3.670 21.890 4.280 ;
        RECT 22.730 3.670 30.630 4.280 ;
        RECT 31.470 3.670 39.830 4.280 ;
        RECT 40.670 3.670 48.570 4.280 ;
        RECT 49.410 3.670 57.770 4.280 ;
        RECT 58.610 3.670 66.510 4.280 ;
        RECT 67.350 3.670 75.710 4.280 ;
        RECT 76.550 3.670 84.450 4.280 ;
        RECT 85.290 3.670 93.650 4.280 ;
        RECT 94.490 3.670 102.390 4.280 ;
        RECT 103.230 3.670 111.590 4.280 ;
        RECT 112.430 3.670 120.330 4.280 ;
        RECT 121.170 3.670 129.530 4.280 ;
        RECT 130.370 3.670 138.270 4.280 ;
        RECT 139.110 3.670 147.470 4.280 ;
        RECT 148.310 3.670 156.670 4.280 ;
        RECT 157.510 3.670 165.410 4.280 ;
        RECT 166.250 3.670 174.610 4.280 ;
        RECT 175.450 3.670 183.350 4.280 ;
        RECT 184.190 3.670 192.550 4.280 ;
        RECT 193.390 3.670 201.290 4.280 ;
        RECT 202.130 3.670 210.490 4.280 ;
        RECT 211.330 3.670 219.230 4.280 ;
        RECT 220.070 3.670 228.430 4.280 ;
        RECT 229.270 3.670 237.170 4.280 ;
        RECT 238.010 3.670 246.370 4.280 ;
        RECT 247.210 3.670 255.110 4.280 ;
        RECT 255.950 3.670 264.310 4.280 ;
        RECT 265.150 3.670 273.050 4.280 ;
        RECT 273.890 3.670 282.250 4.280 ;
        RECT 283.090 3.670 291.450 4.280 ;
        RECT 292.290 3.670 300.190 4.280 ;
        RECT 301.030 3.670 309.390 4.280 ;
        RECT 310.230 3.670 318.130 4.280 ;
        RECT 318.970 3.670 327.330 4.280 ;
        RECT 328.170 3.670 336.070 4.280 ;
        RECT 336.910 3.670 345.270 4.280 ;
        RECT 346.110 3.670 354.010 4.280 ;
        RECT 354.850 3.670 363.210 4.280 ;
        RECT 364.050 3.670 371.950 4.280 ;
        RECT 372.790 3.670 381.150 4.280 ;
        RECT 381.990 3.670 389.890 4.280 ;
        RECT 390.730 3.670 399.090 4.280 ;
        RECT 399.930 3.670 407.830 4.280 ;
        RECT 408.670 3.670 417.030 4.280 ;
        RECT 417.870 3.670 425.770 4.280 ;
        RECT 426.610 3.670 434.970 4.280 ;
        RECT 435.810 3.670 444.170 4.280 ;
        RECT 445.010 3.670 452.910 4.280 ;
        RECT 453.750 3.670 462.110 4.280 ;
        RECT 462.950 3.670 470.850 4.280 ;
        RECT 471.690 3.670 480.050 4.280 ;
        RECT 480.890 3.670 488.790 4.280 ;
        RECT 489.630 3.670 497.990 4.280 ;
        RECT 498.830 3.670 506.730 4.280 ;
        RECT 507.570 3.670 515.930 4.280 ;
        RECT 516.770 3.670 524.670 4.280 ;
        RECT 525.510 3.670 533.870 4.280 ;
        RECT 534.710 3.670 542.610 4.280 ;
        RECT 543.450 3.670 551.810 4.280 ;
        RECT 552.650 3.670 560.550 4.280 ;
        RECT 561.390 3.670 569.750 4.280 ;
        RECT 570.590 3.670 578.950 4.280 ;
        RECT 579.790 3.670 587.690 4.280 ;
        RECT 588.530 3.670 596.890 4.280 ;
        RECT 597.730 3.670 605.630 4.280 ;
        RECT 606.470 3.670 614.830 4.280 ;
        RECT 615.670 3.670 623.570 4.280 ;
        RECT 624.410 3.670 632.770 4.280 ;
        RECT 633.610 3.670 641.510 4.280 ;
        RECT 642.350 3.670 650.710 4.280 ;
        RECT 651.550 3.670 659.450 4.280 ;
        RECT 660.290 3.670 668.650 4.280 ;
        RECT 669.490 3.670 677.390 4.280 ;
        RECT 678.230 3.670 686.590 4.280 ;
        RECT 687.430 3.670 695.330 4.280 ;
        RECT 696.170 3.670 704.530 4.280 ;
        RECT 705.370 3.670 713.270 4.280 ;
        RECT 714.110 3.670 722.470 4.280 ;
        RECT 723.310 3.670 731.670 4.280 ;
        RECT 732.510 3.670 740.410 4.280 ;
        RECT 741.250 3.670 749.610 4.280 ;
        RECT 750.450 3.670 758.350 4.280 ;
        RECT 759.190 3.670 767.550 4.280 ;
        RECT 768.390 3.670 776.290 4.280 ;
        RECT 777.130 3.670 785.490 4.280 ;
        RECT 786.330 3.670 794.230 4.280 ;
        RECT 795.070 3.670 803.430 4.280 ;
        RECT 804.270 3.670 812.170 4.280 ;
        RECT 813.010 3.670 821.370 4.280 ;
        RECT 822.210 3.670 830.110 4.280 ;
        RECT 830.950 3.670 839.310 4.280 ;
        RECT 840.150 3.670 848.050 4.280 ;
        RECT 848.890 3.670 857.250 4.280 ;
        RECT 858.090 3.670 866.450 4.280 ;
        RECT 867.290 3.670 875.190 4.280 ;
        RECT 876.030 3.670 884.390 4.280 ;
        RECT 885.230 3.670 893.130 4.280 ;
        RECT 893.970 3.670 902.330 4.280 ;
        RECT 903.170 3.670 911.070 4.280 ;
        RECT 911.910 3.670 920.270 4.280 ;
        RECT 921.110 3.670 929.010 4.280 ;
        RECT 929.850 3.670 938.210 4.280 ;
        RECT 939.050 3.670 946.950 4.280 ;
        RECT 947.790 3.670 956.150 4.280 ;
        RECT 956.990 3.670 964.890 4.280 ;
        RECT 965.730 3.670 974.090 4.280 ;
        RECT 974.930 3.670 982.830 4.280 ;
        RECT 983.670 3.670 992.030 4.280 ;
        RECT 992.870 3.670 1000.770 4.280 ;
        RECT 1001.610 3.670 1009.970 4.280 ;
        RECT 1010.810 3.670 1019.170 4.280 ;
        RECT 1020.010 3.670 1027.910 4.280 ;
        RECT 1028.750 3.670 1037.110 4.280 ;
        RECT 1037.950 3.670 1045.850 4.280 ;
        RECT 1046.690 3.670 1055.050 4.280 ;
        RECT 1055.890 3.670 1063.790 4.280 ;
        RECT 1064.630 3.670 1072.990 4.280 ;
        RECT 1073.830 3.670 1081.730 4.280 ;
        RECT 1082.570 3.670 1090.930 4.280 ;
        RECT 1091.770 3.670 1099.670 4.280 ;
        RECT 1100.510 3.670 1108.870 4.280 ;
        RECT 1109.710 3.670 1117.610 4.280 ;
        RECT 1118.450 3.670 1126.810 4.280 ;
        RECT 1127.650 3.670 1135.550 4.280 ;
        RECT 1136.390 3.670 1144.750 4.280 ;
        RECT 1145.590 3.670 1149.440 4.280 ;
      LAYER met3 ;
        RECT 4.400 1144.080 1147.175 1144.945 ;
        RECT 3.030 1136.640 1147.175 1144.080 ;
        RECT 4.400 1135.240 1147.175 1136.640 ;
        RECT 3.030 1127.800 1147.175 1135.240 ;
        RECT 4.400 1126.400 1147.175 1127.800 ;
        RECT 3.030 1118.960 1147.175 1126.400 ;
        RECT 4.400 1117.560 1147.175 1118.960 ;
        RECT 3.030 1109.440 1147.175 1117.560 ;
        RECT 4.400 1108.040 1147.175 1109.440 ;
        RECT 3.030 1100.600 1147.175 1108.040 ;
        RECT 4.400 1099.200 1147.175 1100.600 ;
        RECT 3.030 1091.760 1147.175 1099.200 ;
        RECT 4.400 1090.360 1147.175 1091.760 ;
        RECT 3.030 1082.920 1147.175 1090.360 ;
        RECT 4.400 1081.520 1147.175 1082.920 ;
        RECT 3.030 1074.080 1147.175 1081.520 ;
        RECT 4.400 1072.680 1147.175 1074.080 ;
        RECT 3.030 1064.560 1147.175 1072.680 ;
        RECT 4.400 1063.160 1147.175 1064.560 ;
        RECT 3.030 1055.720 1147.175 1063.160 ;
        RECT 4.400 1054.320 1147.175 1055.720 ;
        RECT 3.030 1046.880 1147.175 1054.320 ;
        RECT 4.400 1045.480 1147.175 1046.880 ;
        RECT 3.030 1038.040 1147.175 1045.480 ;
        RECT 4.400 1036.640 1147.175 1038.040 ;
        RECT 3.030 1029.200 1147.175 1036.640 ;
        RECT 4.400 1027.800 1147.175 1029.200 ;
        RECT 3.030 1019.680 1147.175 1027.800 ;
        RECT 4.400 1018.280 1147.175 1019.680 ;
        RECT 3.030 1010.840 1147.175 1018.280 ;
        RECT 4.400 1009.440 1147.175 1010.840 ;
        RECT 3.030 1002.000 1147.175 1009.440 ;
        RECT 4.400 1000.600 1147.175 1002.000 ;
        RECT 3.030 993.160 1147.175 1000.600 ;
        RECT 4.400 991.760 1147.175 993.160 ;
        RECT 3.030 983.640 1147.175 991.760 ;
        RECT 4.400 982.240 1147.175 983.640 ;
        RECT 3.030 974.800 1147.175 982.240 ;
        RECT 4.400 973.400 1147.175 974.800 ;
        RECT 3.030 965.960 1147.175 973.400 ;
        RECT 4.400 964.560 1147.175 965.960 ;
        RECT 3.030 957.120 1147.175 964.560 ;
        RECT 4.400 955.720 1147.175 957.120 ;
        RECT 3.030 948.280 1147.175 955.720 ;
        RECT 4.400 946.880 1147.175 948.280 ;
        RECT 3.030 938.760 1147.175 946.880 ;
        RECT 4.400 937.360 1147.175 938.760 ;
        RECT 3.030 929.920 1147.175 937.360 ;
        RECT 4.400 928.520 1147.175 929.920 ;
        RECT 3.030 921.080 1147.175 928.520 ;
        RECT 4.400 919.680 1147.175 921.080 ;
        RECT 3.030 912.240 1147.175 919.680 ;
        RECT 4.400 910.840 1147.175 912.240 ;
        RECT 3.030 903.400 1147.175 910.840 ;
        RECT 4.400 902.000 1147.175 903.400 ;
        RECT 3.030 893.880 1147.175 902.000 ;
        RECT 4.400 892.480 1147.175 893.880 ;
        RECT 3.030 885.040 1147.175 892.480 ;
        RECT 4.400 883.640 1147.175 885.040 ;
        RECT 3.030 876.200 1147.175 883.640 ;
        RECT 4.400 874.800 1147.175 876.200 ;
        RECT 3.030 867.360 1147.175 874.800 ;
        RECT 4.400 865.960 1147.175 867.360 ;
        RECT 3.030 858.520 1147.175 865.960 ;
        RECT 4.400 857.120 1147.175 858.520 ;
        RECT 3.030 849.000 1147.175 857.120 ;
        RECT 4.400 847.600 1147.175 849.000 ;
        RECT 3.030 840.160 1147.175 847.600 ;
        RECT 4.400 838.760 1147.175 840.160 ;
        RECT 3.030 831.320 1147.175 838.760 ;
        RECT 4.400 829.920 1147.175 831.320 ;
        RECT 3.030 822.480 1147.175 829.920 ;
        RECT 4.400 821.080 1147.175 822.480 ;
        RECT 3.030 812.960 1147.175 821.080 ;
        RECT 4.400 811.560 1147.175 812.960 ;
        RECT 3.030 804.120 1147.175 811.560 ;
        RECT 4.400 802.720 1147.175 804.120 ;
        RECT 3.030 795.280 1147.175 802.720 ;
        RECT 4.400 793.880 1147.175 795.280 ;
        RECT 3.030 786.440 1147.175 793.880 ;
        RECT 4.400 785.040 1147.175 786.440 ;
        RECT 3.030 777.600 1147.175 785.040 ;
        RECT 4.400 776.200 1147.175 777.600 ;
        RECT 3.030 768.080 1147.175 776.200 ;
        RECT 4.400 766.680 1147.175 768.080 ;
        RECT 3.030 759.240 1147.175 766.680 ;
        RECT 4.400 757.840 1147.175 759.240 ;
        RECT 3.030 750.400 1147.175 757.840 ;
        RECT 4.400 749.000 1147.175 750.400 ;
        RECT 3.030 741.560 1147.175 749.000 ;
        RECT 4.400 740.160 1147.175 741.560 ;
        RECT 3.030 732.720 1147.175 740.160 ;
        RECT 4.400 731.320 1147.175 732.720 ;
        RECT 3.030 723.200 1147.175 731.320 ;
        RECT 4.400 721.800 1147.175 723.200 ;
        RECT 3.030 714.360 1147.175 721.800 ;
        RECT 4.400 712.960 1147.175 714.360 ;
        RECT 3.030 705.520 1147.175 712.960 ;
        RECT 4.400 704.120 1147.175 705.520 ;
        RECT 3.030 696.680 1147.175 704.120 ;
        RECT 4.400 695.280 1147.175 696.680 ;
        RECT 3.030 687.840 1147.175 695.280 ;
        RECT 4.400 686.440 1147.175 687.840 ;
        RECT 3.030 678.320 1147.175 686.440 ;
        RECT 4.400 676.920 1147.175 678.320 ;
        RECT 3.030 669.480 1147.175 676.920 ;
        RECT 4.400 668.080 1147.175 669.480 ;
        RECT 3.030 660.640 1147.175 668.080 ;
        RECT 4.400 659.240 1147.175 660.640 ;
        RECT 3.030 651.800 1147.175 659.240 ;
        RECT 4.400 650.400 1147.175 651.800 ;
        RECT 3.030 642.280 1147.175 650.400 ;
        RECT 4.400 640.880 1147.175 642.280 ;
        RECT 3.030 633.440 1147.175 640.880 ;
        RECT 4.400 632.040 1147.175 633.440 ;
        RECT 3.030 624.600 1147.175 632.040 ;
        RECT 4.400 623.200 1147.175 624.600 ;
        RECT 3.030 615.760 1147.175 623.200 ;
        RECT 4.400 614.360 1147.175 615.760 ;
        RECT 3.030 606.920 1147.175 614.360 ;
        RECT 4.400 605.520 1147.175 606.920 ;
        RECT 3.030 597.400 1147.175 605.520 ;
        RECT 4.400 596.000 1147.175 597.400 ;
        RECT 3.030 588.560 1147.175 596.000 ;
        RECT 4.400 587.160 1147.175 588.560 ;
        RECT 3.030 579.720 1147.175 587.160 ;
        RECT 4.400 578.320 1147.175 579.720 ;
        RECT 3.030 570.880 1147.175 578.320 ;
        RECT 4.400 569.480 1147.175 570.880 ;
        RECT 3.030 562.040 1147.175 569.480 ;
        RECT 4.400 560.640 1147.175 562.040 ;
        RECT 3.030 552.520 1147.175 560.640 ;
        RECT 4.400 551.120 1147.175 552.520 ;
        RECT 3.030 543.680 1147.175 551.120 ;
        RECT 4.400 542.280 1147.175 543.680 ;
        RECT 3.030 534.840 1147.175 542.280 ;
        RECT 4.400 533.440 1147.175 534.840 ;
        RECT 3.030 526.000 1147.175 533.440 ;
        RECT 4.400 524.600 1147.175 526.000 ;
        RECT 3.030 517.160 1147.175 524.600 ;
        RECT 4.400 515.760 1147.175 517.160 ;
        RECT 3.030 507.640 1147.175 515.760 ;
        RECT 4.400 506.240 1147.175 507.640 ;
        RECT 3.030 498.800 1147.175 506.240 ;
        RECT 4.400 497.400 1147.175 498.800 ;
        RECT 3.030 489.960 1147.175 497.400 ;
        RECT 4.400 488.560 1147.175 489.960 ;
        RECT 3.030 481.120 1147.175 488.560 ;
        RECT 4.400 479.720 1147.175 481.120 ;
        RECT 3.030 471.600 1147.175 479.720 ;
        RECT 4.400 470.200 1147.175 471.600 ;
        RECT 3.030 462.760 1147.175 470.200 ;
        RECT 4.400 461.360 1147.175 462.760 ;
        RECT 3.030 453.920 1147.175 461.360 ;
        RECT 4.400 452.520 1147.175 453.920 ;
        RECT 3.030 445.080 1147.175 452.520 ;
        RECT 4.400 443.680 1147.175 445.080 ;
        RECT 3.030 436.240 1147.175 443.680 ;
        RECT 4.400 434.840 1147.175 436.240 ;
        RECT 3.030 426.720 1147.175 434.840 ;
        RECT 4.400 425.320 1147.175 426.720 ;
        RECT 3.030 417.880 1147.175 425.320 ;
        RECT 4.400 416.480 1147.175 417.880 ;
        RECT 3.030 409.040 1147.175 416.480 ;
        RECT 4.400 407.640 1147.175 409.040 ;
        RECT 3.030 400.200 1147.175 407.640 ;
        RECT 4.400 398.800 1147.175 400.200 ;
        RECT 3.030 391.360 1147.175 398.800 ;
        RECT 4.400 389.960 1147.175 391.360 ;
        RECT 3.030 381.840 1147.175 389.960 ;
        RECT 4.400 380.440 1147.175 381.840 ;
        RECT 3.030 373.000 1147.175 380.440 ;
        RECT 4.400 371.600 1147.175 373.000 ;
        RECT 3.030 364.160 1147.175 371.600 ;
        RECT 4.400 362.760 1147.175 364.160 ;
        RECT 3.030 355.320 1147.175 362.760 ;
        RECT 4.400 353.920 1147.175 355.320 ;
        RECT 3.030 346.480 1147.175 353.920 ;
        RECT 4.400 345.080 1147.175 346.480 ;
        RECT 3.030 336.960 1147.175 345.080 ;
        RECT 4.400 335.560 1147.175 336.960 ;
        RECT 3.030 328.120 1147.175 335.560 ;
        RECT 4.400 326.720 1147.175 328.120 ;
        RECT 3.030 319.280 1147.175 326.720 ;
        RECT 4.400 317.880 1147.175 319.280 ;
        RECT 3.030 310.440 1147.175 317.880 ;
        RECT 4.400 309.040 1147.175 310.440 ;
        RECT 3.030 300.920 1147.175 309.040 ;
        RECT 4.400 299.520 1147.175 300.920 ;
        RECT 3.030 292.080 1147.175 299.520 ;
        RECT 4.400 290.680 1147.175 292.080 ;
        RECT 3.030 283.240 1147.175 290.680 ;
        RECT 4.400 281.840 1147.175 283.240 ;
        RECT 3.030 274.400 1147.175 281.840 ;
        RECT 4.400 273.000 1147.175 274.400 ;
        RECT 3.030 265.560 1147.175 273.000 ;
        RECT 4.400 264.160 1147.175 265.560 ;
        RECT 3.030 256.040 1147.175 264.160 ;
        RECT 4.400 254.640 1147.175 256.040 ;
        RECT 3.030 247.200 1147.175 254.640 ;
        RECT 4.400 245.800 1147.175 247.200 ;
        RECT 3.030 238.360 1147.175 245.800 ;
        RECT 4.400 236.960 1147.175 238.360 ;
        RECT 3.030 229.520 1147.175 236.960 ;
        RECT 4.400 228.120 1147.175 229.520 ;
        RECT 3.030 220.680 1147.175 228.120 ;
        RECT 4.400 219.280 1147.175 220.680 ;
        RECT 3.030 211.160 1147.175 219.280 ;
        RECT 4.400 209.760 1147.175 211.160 ;
        RECT 3.030 202.320 1147.175 209.760 ;
        RECT 4.400 200.920 1147.175 202.320 ;
        RECT 3.030 193.480 1147.175 200.920 ;
        RECT 4.400 192.080 1147.175 193.480 ;
        RECT 3.030 184.640 1147.175 192.080 ;
        RECT 4.400 183.240 1147.175 184.640 ;
        RECT 3.030 175.800 1147.175 183.240 ;
        RECT 4.400 174.400 1147.175 175.800 ;
        RECT 3.030 166.280 1147.175 174.400 ;
        RECT 4.400 164.880 1147.175 166.280 ;
        RECT 3.030 157.440 1147.175 164.880 ;
        RECT 4.400 156.040 1147.175 157.440 ;
        RECT 3.030 148.600 1147.175 156.040 ;
        RECT 4.400 147.200 1147.175 148.600 ;
        RECT 3.030 139.760 1147.175 147.200 ;
        RECT 4.400 138.360 1147.175 139.760 ;
        RECT 3.030 130.240 1147.175 138.360 ;
        RECT 4.400 128.840 1147.175 130.240 ;
        RECT 3.030 121.400 1147.175 128.840 ;
        RECT 4.400 120.000 1147.175 121.400 ;
        RECT 3.030 112.560 1147.175 120.000 ;
        RECT 4.400 111.160 1147.175 112.560 ;
        RECT 3.030 103.720 1147.175 111.160 ;
        RECT 4.400 102.320 1147.175 103.720 ;
        RECT 3.030 94.880 1147.175 102.320 ;
        RECT 4.400 93.480 1147.175 94.880 ;
        RECT 3.030 85.360 1147.175 93.480 ;
        RECT 4.400 83.960 1147.175 85.360 ;
        RECT 3.030 76.520 1147.175 83.960 ;
        RECT 4.400 75.120 1147.175 76.520 ;
        RECT 3.030 67.680 1147.175 75.120 ;
        RECT 4.400 66.280 1147.175 67.680 ;
        RECT 3.030 58.840 1147.175 66.280 ;
        RECT 4.400 57.440 1147.175 58.840 ;
        RECT 3.030 50.000 1147.175 57.440 ;
        RECT 4.400 48.600 1147.175 50.000 ;
        RECT 3.030 40.480 1147.175 48.600 ;
        RECT 4.400 39.080 1147.175 40.480 ;
        RECT 3.030 31.640 1147.175 39.080 ;
        RECT 4.400 30.240 1147.175 31.640 ;
        RECT 3.030 22.800 1147.175 30.240 ;
        RECT 4.400 21.400 1147.175 22.800 ;
        RECT 3.030 13.960 1147.175 21.400 ;
        RECT 4.400 12.560 1147.175 13.960 ;
        RECT 3.030 5.120 1147.175 12.560 ;
        RECT 4.400 4.255 1147.175 5.120 ;
      LAYER met4 ;
        RECT 3.055 1137.600 1135.905 1138.145 ;
        RECT 3.055 10.240 8.570 1137.600 ;
        RECT 12.470 10.240 98.570 1137.600 ;
        RECT 102.470 10.240 188.570 1137.600 ;
        RECT 192.470 10.240 278.570 1137.600 ;
        RECT 282.470 10.240 368.570 1137.600 ;
        RECT 372.470 10.240 458.570 1137.600 ;
        RECT 462.470 10.240 548.570 1137.600 ;
        RECT 552.470 10.240 638.570 1137.600 ;
        RECT 642.470 10.240 728.570 1137.600 ;
        RECT 732.470 10.240 818.570 1137.600 ;
        RECT 822.470 10.240 908.570 1137.600 ;
        RECT 912.470 10.240 998.570 1137.600 ;
        RECT 1002.470 10.240 1088.570 1137.600 ;
        RECT 1092.470 10.240 1135.905 1137.600 ;
        RECT 3.055 8.335 1135.905 10.240 ;
  END
END Microwatt_FP_DFFRFile
END LIBRARY

