VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM512
  CLASS BLOCK ;
  FOREIGN RAM512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1594.820 BY 987.360 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 520.920 1594.820 521.520 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 575.320 1594.820 575.920 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 630.400 1594.820 631.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 685.480 1594.820 686.080 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 739.880 1594.820 740.480 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 794.960 1594.820 795.560 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 850.040 1594.820 850.640 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 904.440 1594.820 905.040 ;
    END
  END A0[7]
  PIN A0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 959.520 1594.820 960.120 ;
    END
  END A0[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 2.000 494.320 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 0.000 710.150 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 0.000 934.630 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 0.000 959.470 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 0.000 984.310 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 0.000 1009.150 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 0.000 1108.970 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.370 0.000 1158.650 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 0.000 1258.470 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 0.000 1308.150 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 0.000 1358.290 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 0.000 1383.130 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 0.000 1407.970 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.530 0.000 1432.810 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 0.000 1457.650 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.670 0.000 1482.950 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 0.000 1507.790 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.350 0.000 1532.630 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 0.000 1557.470 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.030 0.000 1582.310 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 985.360 12.790 987.360 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 985.360 261.650 987.360 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 985.360 286.490 987.360 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 985.360 311.790 987.360 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 985.360 336.630 987.360 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 985.360 361.470 987.360 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 985.360 386.310 987.360 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 985.360 411.150 987.360 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 985.360 435.990 987.360 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 985.360 461.290 987.360 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 985.360 486.130 987.360 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 985.360 37.630 987.360 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 985.360 510.970 987.360 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 985.360 535.810 987.360 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 985.360 560.650 987.360 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 985.360 585.490 987.360 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 985.360 610.790 987.360 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 985.360 635.630 987.360 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 985.360 660.470 987.360 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 985.360 685.310 987.360 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 985.360 710.150 987.360 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 985.360 734.990 987.360 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 985.360 62.470 987.360 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 985.360 760.290 987.360 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 985.360 785.130 987.360 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 985.360 809.970 987.360 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 985.360 834.810 987.360 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 985.360 859.650 987.360 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 985.360 884.950 987.360 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 985.360 909.790 987.360 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 985.360 934.630 987.360 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 985.360 959.470 987.360 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 985.360 984.310 987.360 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 985.360 87.310 987.360 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 985.360 1009.150 987.360 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 985.360 1034.450 987.360 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 985.360 1059.290 987.360 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 985.360 1084.130 987.360 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 985.360 1108.970 987.360 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 985.360 1133.810 987.360 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.370 985.360 1158.650 987.360 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 985.360 1183.950 987.360 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 985.360 1208.790 987.360 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 985.360 1233.630 987.360 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 985.360 112.150 987.360 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 985.360 1258.470 987.360 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 985.360 1283.310 987.360 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 985.360 1308.150 987.360 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 985.360 1333.450 987.360 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 985.360 1358.290 987.360 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 985.360 1383.130 987.360 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 985.360 1407.970 987.360 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.530 985.360 1432.810 987.360 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 985.360 1457.650 987.360 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.670 985.360 1482.950 987.360 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 985.360 136.990 987.360 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 985.360 1507.790 987.360 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.350 985.360 1532.630 987.360 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 985.360 1557.470 987.360 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.030 985.360 1582.310 987.360 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 985.360 162.290 987.360 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 985.360 187.130 987.360 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 985.360 211.970 987.360 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 985.360 236.810 987.360 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 27.240 1594.820 27.840 ;
    END
  END EN0
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 113.690 100.400 116.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.690 100.400 296.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.690 100.400 476.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.690 100.400 656.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 833.690 100.400 836.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.690 100.400 1016.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.690 100.400 1196.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.690 100.400 1376.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1553.690 100.400 1556.790 886.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.690 100.400 26.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.690 100.400 206.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.690 100.400 386.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.690 100.400 566.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.690 100.400 746.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.690 100.400 926.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.690 100.400 1106.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.690 100.400 1286.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.690 100.400 1466.790 886.960 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 81.640 1594.820 82.240 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 136.720 1594.820 137.320 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 191.800 1594.820 192.400 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 246.200 1594.820 246.800 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 301.280 1594.820 301.880 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 356.360 1594.820 356.960 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 410.760 1594.820 411.360 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1592.820 465.840 1594.820 466.440 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 20.240 100.555 1574.580 886.805 ;
      LAYER met1 ;
        RECT 1.450 0.040 1593.370 987.320 ;
      LAYER met2 ;
        RECT 1.480 985.080 12.230 987.350 ;
        RECT 13.070 985.080 37.070 987.350 ;
        RECT 37.910 985.080 61.910 987.350 ;
        RECT 62.750 985.080 86.750 987.350 ;
        RECT 87.590 985.080 111.590 987.350 ;
        RECT 112.430 985.080 136.430 987.350 ;
        RECT 137.270 985.080 161.730 987.350 ;
        RECT 162.570 985.080 186.570 987.350 ;
        RECT 187.410 985.080 211.410 987.350 ;
        RECT 212.250 985.080 236.250 987.350 ;
        RECT 237.090 985.080 261.090 987.350 ;
        RECT 261.930 985.080 285.930 987.350 ;
        RECT 286.770 985.080 311.230 987.350 ;
        RECT 312.070 985.080 336.070 987.350 ;
        RECT 336.910 985.080 360.910 987.350 ;
        RECT 361.750 985.080 385.750 987.350 ;
        RECT 386.590 985.080 410.590 987.350 ;
        RECT 411.430 985.080 435.430 987.350 ;
        RECT 436.270 985.080 460.730 987.350 ;
        RECT 461.570 985.080 485.570 987.350 ;
        RECT 486.410 985.080 510.410 987.350 ;
        RECT 511.250 985.080 535.250 987.350 ;
        RECT 536.090 985.080 560.090 987.350 ;
        RECT 560.930 985.080 584.930 987.350 ;
        RECT 585.770 985.080 610.230 987.350 ;
        RECT 611.070 985.080 635.070 987.350 ;
        RECT 635.910 985.080 659.910 987.350 ;
        RECT 660.750 985.080 684.750 987.350 ;
        RECT 685.590 985.080 709.590 987.350 ;
        RECT 710.430 985.080 734.430 987.350 ;
        RECT 735.270 985.080 759.730 987.350 ;
        RECT 760.570 985.080 784.570 987.350 ;
        RECT 785.410 985.080 809.410 987.350 ;
        RECT 810.250 985.080 834.250 987.350 ;
        RECT 835.090 985.080 859.090 987.350 ;
        RECT 859.930 985.080 884.390 987.350 ;
        RECT 885.230 985.080 909.230 987.350 ;
        RECT 910.070 985.080 934.070 987.350 ;
        RECT 934.910 985.080 958.910 987.350 ;
        RECT 959.750 985.080 983.750 987.350 ;
        RECT 984.590 985.080 1008.590 987.350 ;
        RECT 1009.430 985.080 1033.890 987.350 ;
        RECT 1034.730 985.080 1058.730 987.350 ;
        RECT 1059.570 985.080 1083.570 987.350 ;
        RECT 1084.410 985.080 1108.410 987.350 ;
        RECT 1109.250 985.080 1133.250 987.350 ;
        RECT 1134.090 985.080 1158.090 987.350 ;
        RECT 1158.930 985.080 1183.390 987.350 ;
        RECT 1184.230 985.080 1208.230 987.350 ;
        RECT 1209.070 985.080 1233.070 987.350 ;
        RECT 1233.910 985.080 1257.910 987.350 ;
        RECT 1258.750 985.080 1282.750 987.350 ;
        RECT 1283.590 985.080 1307.590 987.350 ;
        RECT 1308.430 985.080 1332.890 987.350 ;
        RECT 1333.730 985.080 1357.730 987.350 ;
        RECT 1358.570 985.080 1382.570 987.350 ;
        RECT 1383.410 985.080 1407.410 987.350 ;
        RECT 1408.250 985.080 1432.250 987.350 ;
        RECT 1433.090 985.080 1457.090 987.350 ;
        RECT 1457.930 985.080 1482.390 987.350 ;
        RECT 1483.230 985.080 1507.230 987.350 ;
        RECT 1508.070 985.080 1532.070 987.350 ;
        RECT 1532.910 985.080 1556.910 987.350 ;
        RECT 1557.750 985.080 1581.750 987.350 ;
        RECT 1582.590 985.080 1593.340 987.350 ;
        RECT 1.480 2.280 1593.340 985.080 ;
        RECT 1.480 0.010 12.230 2.280 ;
        RECT 13.070 0.010 37.070 2.280 ;
        RECT 37.910 0.010 61.910 2.280 ;
        RECT 62.750 0.010 86.750 2.280 ;
        RECT 87.590 0.010 111.590 2.280 ;
        RECT 112.430 0.010 136.430 2.280 ;
        RECT 137.270 0.010 161.730 2.280 ;
        RECT 162.570 0.010 186.570 2.280 ;
        RECT 187.410 0.010 211.410 2.280 ;
        RECT 212.250 0.010 236.250 2.280 ;
        RECT 237.090 0.010 261.090 2.280 ;
        RECT 261.930 0.010 285.930 2.280 ;
        RECT 286.770 0.010 311.230 2.280 ;
        RECT 312.070 0.010 336.070 2.280 ;
        RECT 336.910 0.010 360.910 2.280 ;
        RECT 361.750 0.010 385.750 2.280 ;
        RECT 386.590 0.010 410.590 2.280 ;
        RECT 411.430 0.010 435.430 2.280 ;
        RECT 436.270 0.010 460.730 2.280 ;
        RECT 461.570 0.010 485.570 2.280 ;
        RECT 486.410 0.010 510.410 2.280 ;
        RECT 511.250 0.010 535.250 2.280 ;
        RECT 536.090 0.010 560.090 2.280 ;
        RECT 560.930 0.010 584.930 2.280 ;
        RECT 585.770 0.010 610.230 2.280 ;
        RECT 611.070 0.010 635.070 2.280 ;
        RECT 635.910 0.010 659.910 2.280 ;
        RECT 660.750 0.010 684.750 2.280 ;
        RECT 685.590 0.010 709.590 2.280 ;
        RECT 710.430 0.010 734.430 2.280 ;
        RECT 735.270 0.010 759.730 2.280 ;
        RECT 760.570 0.010 784.570 2.280 ;
        RECT 785.410 0.010 809.410 2.280 ;
        RECT 810.250 0.010 834.250 2.280 ;
        RECT 835.090 0.010 859.090 2.280 ;
        RECT 859.930 0.010 884.390 2.280 ;
        RECT 885.230 0.010 909.230 2.280 ;
        RECT 910.070 0.010 934.070 2.280 ;
        RECT 934.910 0.010 958.910 2.280 ;
        RECT 959.750 0.010 983.750 2.280 ;
        RECT 984.590 0.010 1008.590 2.280 ;
        RECT 1009.430 0.010 1033.890 2.280 ;
        RECT 1034.730 0.010 1058.730 2.280 ;
        RECT 1059.570 0.010 1083.570 2.280 ;
        RECT 1084.410 0.010 1108.410 2.280 ;
        RECT 1109.250 0.010 1133.250 2.280 ;
        RECT 1134.090 0.010 1158.090 2.280 ;
        RECT 1158.930 0.010 1183.390 2.280 ;
        RECT 1184.230 0.010 1208.230 2.280 ;
        RECT 1209.070 0.010 1233.070 2.280 ;
        RECT 1233.910 0.010 1257.910 2.280 ;
        RECT 1258.750 0.010 1282.750 2.280 ;
        RECT 1283.590 0.010 1307.590 2.280 ;
        RECT 1308.430 0.010 1332.890 2.280 ;
        RECT 1333.730 0.010 1357.730 2.280 ;
        RECT 1358.570 0.010 1382.570 2.280 ;
        RECT 1383.410 0.010 1407.410 2.280 ;
        RECT 1408.250 0.010 1432.250 2.280 ;
        RECT 1433.090 0.010 1457.090 2.280 ;
        RECT 1457.930 0.010 1482.390 2.280 ;
        RECT 1483.230 0.010 1507.230 2.280 ;
        RECT 1508.070 0.010 1532.070 2.280 ;
        RECT 1532.910 0.010 1556.910 2.280 ;
        RECT 1557.750 0.010 1581.750 2.280 ;
        RECT 1582.590 0.010 1593.340 2.280 ;
      LAYER met3 ;
        RECT 2.000 960.520 1592.820 987.185 ;
        RECT 2.000 959.120 1592.420 960.520 ;
        RECT 2.000 905.440 1592.820 959.120 ;
        RECT 2.000 904.040 1592.420 905.440 ;
        RECT 2.000 851.040 1592.820 904.040 ;
        RECT 2.000 849.640 1592.420 851.040 ;
        RECT 2.000 795.960 1592.820 849.640 ;
        RECT 2.000 794.560 1592.420 795.960 ;
        RECT 2.000 740.880 1592.820 794.560 ;
        RECT 2.000 739.480 1592.420 740.880 ;
        RECT 2.000 686.480 1592.820 739.480 ;
        RECT 2.000 685.080 1592.420 686.480 ;
        RECT 2.000 631.400 1592.820 685.080 ;
        RECT 2.000 630.000 1592.420 631.400 ;
        RECT 2.000 576.320 1592.820 630.000 ;
        RECT 2.000 574.920 1592.420 576.320 ;
        RECT 2.000 521.920 1592.820 574.920 ;
        RECT 2.000 520.520 1592.420 521.920 ;
        RECT 2.000 494.720 1592.820 520.520 ;
        RECT 2.400 493.320 1592.820 494.720 ;
        RECT 2.000 466.840 1592.820 493.320 ;
        RECT 2.000 465.440 1592.420 466.840 ;
        RECT 2.000 411.760 1592.820 465.440 ;
        RECT 2.000 410.360 1592.420 411.760 ;
        RECT 2.000 357.360 1592.820 410.360 ;
        RECT 2.000 355.960 1592.420 357.360 ;
        RECT 2.000 302.280 1592.820 355.960 ;
        RECT 2.000 300.880 1592.420 302.280 ;
        RECT 2.000 247.200 1592.820 300.880 ;
        RECT 2.000 245.800 1592.420 247.200 ;
        RECT 2.000 192.800 1592.820 245.800 ;
        RECT 2.000 191.400 1592.420 192.800 ;
        RECT 2.000 137.720 1592.820 191.400 ;
        RECT 2.000 136.320 1592.420 137.720 ;
        RECT 2.000 82.640 1592.820 136.320 ;
        RECT 2.000 81.240 1592.420 82.640 ;
        RECT 2.000 28.240 1592.820 81.240 ;
        RECT 2.000 26.840 1592.420 28.240 ;
        RECT 2.000 0.175 1592.820 26.840 ;
      LAYER met4 ;
        RECT 4.895 887.360 1566.465 987.185 ;
        RECT 4.895 100.000 23.290 887.360 ;
        RECT 27.190 100.000 113.290 887.360 ;
        RECT 117.190 100.000 203.290 887.360 ;
        RECT 207.190 100.000 293.290 887.360 ;
        RECT 297.190 100.000 383.290 887.360 ;
        RECT 387.190 100.000 473.290 887.360 ;
        RECT 477.190 100.000 563.290 887.360 ;
        RECT 567.190 100.000 653.290 887.360 ;
        RECT 657.190 100.000 743.290 887.360 ;
        RECT 747.190 100.000 833.290 887.360 ;
        RECT 837.190 100.000 923.290 887.360 ;
        RECT 927.190 100.000 1013.290 887.360 ;
        RECT 1017.190 100.000 1103.290 887.360 ;
        RECT 1107.190 100.000 1193.290 887.360 ;
        RECT 1197.190 100.000 1283.290 887.360 ;
        RECT 1287.190 100.000 1373.290 887.360 ;
        RECT 1377.190 100.000 1463.290 887.360 ;
        RECT 1467.190 100.000 1553.290 887.360 ;
        RECT 1557.190 100.000 1566.465 887.360 ;
        RECT 4.895 0.855 1566.465 100.000 ;
  END
END RAM512
END LIBRARY

